
module mul_DW_mult_uns_1 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n302, n303, n304, n305, n306, n307, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n817, n820, n823, n826, n829, n832, n835, n838, n841, n844,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311;

  XOR2X1TF U226 ( .A(n227), .B(n226), .Y(product[63]) );
  XOR2X1TF U227 ( .A(n2289), .B(n291), .Y(n226) );
  CMPR32X2TF U228 ( .A(n292), .B(n293), .C(n228), .CO(n227), .S(product[62])
         );
  CMPR32X2TF U229 ( .A(n295), .B(n294), .C(n229), .CO(n228), .S(product[61])
         );
  CMPR32X2TF U230 ( .A(n299), .B(n296), .C(n230), .CO(n229), .S(product[60])
         );
  CMPR32X2TF U231 ( .A(n300), .B(n302), .C(n231), .CO(n230), .S(product[59])
         );
  CMPR32X2TF U232 ( .A(n303), .B(n305), .C(n232), .CO(n231), .S(product[58])
         );
  CMPR32X2TF U233 ( .A(n306), .B(n310), .C(n233), .CO(n232), .S(product[57])
         );
  CMPR32X2TF U234 ( .A(n311), .B(n314), .C(n234), .CO(n233), .S(product[56])
         );
  CMPR32X2TF U235 ( .A(n315), .B(n318), .C(n235), .CO(n234), .S(product[55])
         );
  CMPR32X2TF U236 ( .A(n319), .B(n325), .C(n236), .CO(n235), .S(product[54])
         );
  CMPR32X2TF U237 ( .A(n326), .B(n331), .C(n237), .CO(n236), .S(product[53])
         );
  CMPR32X2TF U238 ( .A(n332), .B(n336), .C(n238), .CO(n237), .S(product[52])
         );
  CMPR32X2TF U239 ( .A(n337), .B(n344), .C(n239), .CO(n238), .S(product[51])
         );
  CMPR32X2TF U240 ( .A(n345), .B(n351), .C(n240), .CO(n239), .S(product[50])
         );
  CMPR32X2TF U241 ( .A(n352), .B(n359), .C(n241), .CO(n240), .S(product[49])
         );
  CMPR32X2TF U242 ( .A(n360), .B(n369), .C(n242), .CO(n241), .S(product[48])
         );
  CMPR32X2TF U243 ( .A(n370), .B(n378), .C(n243), .CO(n242), .S(product[47])
         );
  CMPR32X2TF U244 ( .A(n379), .B(n386), .C(n244), .CO(n243), .S(product[46])
         );
  CMPR32X2TF U245 ( .A(n387), .B(n397), .C(n245), .CO(n244), .S(product[45])
         );
  CMPR32X2TF U246 ( .A(n398), .B(n407), .C(n246), .CO(n245), .S(product[44])
         );
  CMPR32X2TF U247 ( .A(n408), .B(n418), .C(n247), .CO(n246), .S(product[43])
         );
  CMPR32X2TF U248 ( .A(n419), .B(n431), .C(n248), .CO(n247), .S(product[42])
         );
  CMPR32X2TF U249 ( .A(n432), .B(n443), .C(n249), .CO(n248), .S(product[41])
         );
  CMPR32X2TF U250 ( .A(n444), .B(n454), .C(n250), .CO(n249), .S(product[40])
         );
  CMPR32X2TF U251 ( .A(n455), .B(n468), .C(n251), .CO(n250), .S(product[39])
         );
  CMPR32X2TF U252 ( .A(n469), .B(n481), .C(n252), .CO(n251), .S(product[38])
         );
  CMPR32X2TF U253 ( .A(n482), .B(n495), .C(n253), .CO(n252), .S(product[37])
         );
  CMPR32X2TF U254 ( .A(n496), .B(n509), .C(n254), .CO(n253), .S(product[36])
         );
  CMPR32X2TF U255 ( .A(n510), .B(n1224), .C(n255), .CO(n254), .S(product[35])
         );
  CMPR32X2TF U256 ( .A(n524), .B(n537), .C(n256), .CO(n255), .S(product[34])
         );
  CMPR32X2TF U257 ( .A(n538), .B(n1258), .C(n257), .CO(n256), .S(product[33])
         );
  CMPR32X2TF U258 ( .A(n1259), .B(n552), .C(n258), .CO(n257), .S(product[32])
         );
  CMPR32X2TF U259 ( .A(n1260), .B(n566), .C(n259), .CO(n258), .S(product[31])
         );
  CMPR32X2TF U260 ( .A(n1261), .B(n580), .C(n260), .CO(n259), .S(product[30])
         );
  CMPR32X2TF U261 ( .A(n1262), .B(n594), .C(n261), .CO(n260), .S(product[29])
         );
  CMPR32X2TF U262 ( .A(n1263), .B(n608), .C(n262), .CO(n261), .S(product[28])
         );
  CMPR32X2TF U263 ( .A(n1264), .B(n622), .C(n263), .CO(n262), .S(product[27])
         );
  CMPR32X2TF U264 ( .A(n1265), .B(n636), .C(n264), .CO(n263), .S(product[26])
         );
  CMPR32X2TF U265 ( .A(n1266), .B(n649), .C(n265), .CO(n264), .S(product[25])
         );
  CMPR32X2TF U266 ( .A(n1267), .B(n662), .C(n266), .CO(n265), .S(product[24])
         );
  CMPR32X2TF U267 ( .A(n1268), .B(n675), .C(n267), .CO(n266), .S(product[23])
         );
  CMPR32X2TF U268 ( .A(n1269), .B(n686), .C(n268), .CO(n267), .S(product[22])
         );
  CMPR32X2TF U269 ( .A(n1270), .B(n697), .C(n269), .CO(n268), .S(product[21])
         );
  CMPR32X2TF U270 ( .A(n1271), .B(n708), .C(n270), .CO(n269), .S(product[20])
         );
  CMPR32X2TF U271 ( .A(n1272), .B(n718), .C(n271), .CO(n270), .S(product[19])
         );
  CMPR32X2TF U272 ( .A(n1273), .B(n728), .C(n272), .CO(n271), .S(product[18])
         );
  CMPR32X2TF U273 ( .A(n1274), .B(n738), .C(n273), .CO(n272), .S(product[17])
         );
  CMPR32X2TF U274 ( .A(n1275), .B(n746), .C(n274), .CO(n273), .S(product[16])
         );
  CMPR32X2TF U275 ( .A(n1276), .B(n754), .C(n275), .CO(n274), .S(product[15])
         );
  CMPR32X2TF U276 ( .A(n1277), .B(n762), .C(n276), .CO(n275), .S(product[14])
         );
  CMPR32X2TF U277 ( .A(n1278), .B(n769), .C(n277), .CO(n276), .S(product[13])
         );
  CMPR32X2TF U278 ( .A(n1279), .B(n776), .C(n278), .CO(n277), .S(product[12])
         );
  CMPR32X2TF U279 ( .A(n1280), .B(n783), .C(n279), .CO(n278), .S(product[11])
         );
  CMPR32X2TF U280 ( .A(n1281), .B(n788), .C(n280), .CO(n279), .S(product[10])
         );
  CMPR32X2TF U281 ( .A(n1282), .B(n793), .C(n281), .CO(n280), .S(product[9])
         );
  CMPR32X2TF U282 ( .A(n1283), .B(n797), .C(n282), .CO(n281), .S(product[8])
         );
  CMPR32X2TF U283 ( .A(n1284), .B(n801), .C(n283), .CO(n282), .S(product[7])
         );
  CMPR32X2TF U284 ( .A(n1285), .B(n805), .C(n284), .CO(n283), .S(product[6])
         );
  CMPR32X2TF U285 ( .A(n1286), .B(n809), .C(n285), .CO(n284), .S(product[5])
         );
  CMPR32X2TF U286 ( .A(n1287), .B(n811), .C(n286), .CO(n285), .S(product[4])
         );
  CMPR32X2TF U287 ( .A(n1288), .B(n813), .C(n287), .CO(n286), .S(product[3])
         );
  ADDHXLTF U288 ( .A(n1289), .B(n288), .CO(n287), .S(product[2]) );
  ADDHXLTF U289 ( .A(n1290), .B(n289), .CO(n288), .S(product[1]) );
  ADDHXLTF U290 ( .A(n7), .B(n1291), .CO(n289), .S(product[0]) );
  INVX2TF U292 ( .A(n291), .Y(n292) );
  CMPR32X2TF U293 ( .A(n297), .B(n942), .C(n913), .CO(n293), .S(n294) );
  CMPR32X2TF U294 ( .A(n914), .B(n298), .C(n943), .CO(n295), .S(n296) );
  INVX2TF U295 ( .A(n297), .Y(n298) );
  CMPR32X2TF U296 ( .A(n298), .B(n915), .C(n944), .CO(n299), .S(n300) );
  CMPR42X1TF U298 ( .A(n977), .B(n307), .C(n916), .D(n304), .ICI(n945), .S(
        n303), .ICO(n297), .CO(n302) );
  CMPR42X1TF U299 ( .A(n312), .B(n917), .C(n309), .D(n946), .ICI(n978), .S(
        n306), .ICO(n304), .CO(n305) );
  CMPR42X1TF U301 ( .A(n918), .B(n312), .C(n947), .D(n313), .ICI(n979), .S(
        n311), .ICO(n309), .CO(n310) );
  INVX2TF U302 ( .A(n307), .Y(n312) );
  CMPR42X1TF U303 ( .A(n316), .B(n320), .C(n948), .D(n317), .ICI(n980), .S(
        n315), .ICO(n313), .CO(n314) );
  CMPR32X2TF U304 ( .A(n322), .B(n1012), .C(n919), .CO(n307), .S(n316) );
  CMPR42X1TF U305 ( .A(n949), .B(n321), .C(n324), .D(n981), .ICI(n1013), .S(
        n319), .ICO(n317), .CO(n318) );
  CMPR32X2TF U306 ( .A(n920), .B(n323), .C(n327), .CO(n320), .S(n321) );
  INVX2TF U307 ( .A(n322), .Y(n323) );
  CMPR42X1TF U308 ( .A(n333), .B(n328), .C(n330), .D(n982), .ICI(n1014), .S(
        n326), .ICO(n324), .CO(n325) );
  CMPR32X2TF U309 ( .A(n323), .B(n921), .C(n950), .CO(n327), .S(n328) );
  CMPR42X1TF U311 ( .A(n334), .B(n339), .C(n983), .D(n335), .ICI(n1015), .S(
        n332), .ICO(n330), .CO(n331) );
  CMPR42X1TF U312 ( .A(n1047), .B(n341), .C(n922), .D(n338), .ICI(n951), .S(
        n334), .ICO(n322), .CO(n333) );
  CMPR42X1TF U313 ( .A(n984), .B(n340), .C(n343), .D(n1016), .ICI(n1048), .S(
        n337), .ICO(n335), .CO(n336) );
  CMPR42X1TF U314 ( .A(n349), .B(n923), .C(n346), .D(n952), .ICI(n347), .S(
        n340), .ICO(n338), .CO(n339) );
  CMPR42X1TF U316 ( .A(n354), .B(n348), .C(n350), .D(n1017), .ICI(n1049), .S(
        n345), .ICO(n343), .CO(n344) );
  CMPR42X1TF U317 ( .A(n356), .B(n349), .C(n953), .D(n353), .ICI(n985), .S(
        n348), .ICO(n346), .CO(n347) );
  INVX2TF U318 ( .A(n341), .Y(n349) );
  CMPR42X1TF U319 ( .A(n355), .B(n362), .C(n1018), .D(n358), .ICI(n1050), .S(
        n352), .ICO(n350), .CO(n351) );
  CMPR42X1TF U320 ( .A(n357), .B(n364), .C(n954), .D(n361), .ICI(n986), .S(
        n355), .ICO(n353), .CO(n354) );
  CMPR32X2TF U321 ( .A(n366), .B(n1082), .C(n924), .CO(n356), .S(n357) );
  CMPR42X1TF U322 ( .A(n1019), .B(n363), .C(n368), .D(n1051), .ICI(n1083), .S(
        n360), .ICO(n358), .CO(n359) );
  CMPR42X1TF U323 ( .A(n374), .B(n365), .C(n371), .D(n987), .ICI(n372), .S(
        n363), .ICO(n361), .CO(n362) );
  CMPR32X2TF U324 ( .A(n925), .B(n367), .C(n955), .CO(n364), .S(n365) );
  INVX2TF U325 ( .A(n366), .Y(n367) );
  CMPR42X1TF U326 ( .A(n381), .B(n373), .C(n377), .D(n1052), .ICI(n1084), .S(
        n370), .ICO(n368), .CO(n369) );
  CMPR42X1TF U327 ( .A(n383), .B(n375), .C(n380), .D(n988), .ICI(n1020), .S(
        n373), .ICO(n371), .CO(n372) );
  CMPR32X2TF U328 ( .A(n367), .B(n926), .C(n956), .CO(n374), .S(n375) );
  CMPR42X1TF U330 ( .A(n382), .B(n389), .C(n1053), .D(n385), .ICI(n1085), .S(
        n379), .ICO(n377), .CO(n378) );
  CMPR42X1TF U331 ( .A(n384), .B(n392), .C(n989), .D(n388), .ICI(n1021), .S(
        n382), .ICO(n380), .CO(n381) );
  CMPR42X1TF U332 ( .A(n1117), .B(n394), .C(n927), .D(n391), .ICI(n957), .S(
        n384), .ICO(n366), .CO(n383) );
  CMPR42X1TF U333 ( .A(n1054), .B(n390), .C(n396), .D(n1086), .ICI(n1118), .S(
        n387), .ICO(n385), .CO(n386) );
  CMPR42X1TF U334 ( .A(n990), .B(n393), .C(n399), .D(n1022), .ICI(n400), .S(
        n390), .ICO(n388), .CO(n389) );
  CMPR42X1TF U335 ( .A(n405), .B(n928), .C(n402), .D(n958), .ICI(n403), .S(
        n393), .ICO(n391), .CO(n392) );
  CMPR42X1TF U337 ( .A(n410), .B(n401), .C(n406), .D(n1087), .ICI(n1119), .S(
        n398), .ICO(n396), .CO(n397) );
  CMPR42X1TF U338 ( .A(n413), .B(n404), .C(n409), .D(n1023), .ICI(n1055), .S(
        n401), .ICO(n399), .CO(n400) );
  CMPR42X1TF U339 ( .A(n415), .B(n405), .C(n959), .D(n412), .ICI(n991), .S(
        n404), .ICO(n402), .CO(n403) );
  INVX2TF U340 ( .A(n394), .Y(n405) );
  CMPR42X1TF U341 ( .A(n411), .B(n421), .C(n1088), .D(n417), .ICI(n1120), .S(
        n408), .ICO(n406), .CO(n407) );
  CMPR42X1TF U342 ( .A(n414), .B(n424), .C(n1024), .D(n420), .ICI(n1056), .S(
        n411), .ICO(n409), .CO(n410) );
  CMPR42X1TF U343 ( .A(n416), .B(n960), .C(n426), .D(n423), .ICI(n992), .S(
        n414), .ICO(n412), .CO(n413) );
  CMPR32X2TF U344 ( .A(n428), .B(n1152), .C(n929), .CO(n415), .S(n416) );
  CMPR42X1TF U345 ( .A(n1089), .B(n422), .C(n430), .D(n1121), .ICI(n1153), .S(
        n419), .ICO(n417), .CO(n418) );
  CMPR42X1TF U346 ( .A(n1025), .B(n425), .C(n433), .D(n1057), .ICI(n434), .S(
        n422), .ICO(n420), .CO(n421) );
  CMPR42X1TF U347 ( .A(n439), .B(n427), .C(n436), .D(n993), .ICI(n437), .S(
        n425), .ICO(n423), .CO(n424) );
  CMPR32X2TF U348 ( .A(n930), .B(n429), .C(n961), .CO(n426), .S(n427) );
  INVX2TF U349 ( .A(n428), .Y(n429) );
  CMPR42X1TF U350 ( .A(n446), .B(n435), .C(n442), .D(n1122), .ICI(n1154), .S(
        n432), .ICO(n430), .CO(n431) );
  CMPR42X1TF U351 ( .A(n449), .B(n438), .C(n445), .D(n1058), .ICI(n1090), .S(
        n435), .ICO(n433), .CO(n434) );
  CMPR42X1TF U352 ( .A(n451), .B(n440), .C(n448), .D(n994), .ICI(n1026), .S(
        n438), .ICO(n436), .CO(n437) );
  CMPR32X2TF U353 ( .A(n429), .B(n931), .C(n962), .CO(n439), .S(n440) );
  CMPR42X1TF U355 ( .A(n447), .B(n457), .C(n1123), .D(n453), .ICI(n1155), .S(
        n444), .ICO(n442), .CO(n443) );
  CMPR42X1TF U356 ( .A(n450), .B(n460), .C(n1059), .D(n456), .ICI(n1091), .S(
        n447), .ICO(n445), .CO(n446) );
  CMPR42X1TF U357 ( .A(n452), .B(n463), .C(n995), .D(n459), .ICI(n1027), .S(
        n450), .ICO(n448), .CO(n449) );
  CMPR42X1TF U358 ( .A(n1187), .B(n465), .C(n932), .D(n462), .ICI(n963), .S(
        n452), .ICO(n428), .CO(n451) );
  CMPR42X1TF U359 ( .A(n1124), .B(n458), .C(n467), .D(n1156), .ICI(n1188), .S(
        n455), .ICO(n453), .CO(n454) );
  CMPR42X1TF U360 ( .A(n1060), .B(n461), .C(n470), .D(n1092), .ICI(n471), .S(
        n458), .ICO(n456), .CO(n457) );
  CMPR42X1TF U361 ( .A(n996), .B(n464), .C(n473), .D(n1028), .ICI(n474), .S(
        n461), .ICO(n459), .CO(n460) );
  CMPR42X1TF U362 ( .A(n479), .B(n933), .C(n476), .D(n964), .ICI(n477), .S(
        n464), .ICO(n462), .CO(n463) );
  CMPR42X1TF U364 ( .A(n484), .B(n472), .C(n480), .D(n1157), .ICI(n1189), .S(
        n469), .ICO(n467), .CO(n468) );
  CMPR42X1TF U365 ( .A(n487), .B(n475), .C(n483), .D(n1093), .ICI(n1125), .S(
        n472), .ICO(n470), .CO(n471) );
  CMPR42X1TF U366 ( .A(n490), .B(n478), .C(n486), .D(n1029), .ICI(n1061), .S(
        n475), .ICO(n473), .CO(n474) );
  CMPR42X1TF U367 ( .A(n492), .B(n479), .C(n965), .D(n489), .ICI(n997), .S(
        n478), .ICO(n476), .CO(n477) );
  INVX2TF U368 ( .A(n465), .Y(n479) );
  CMPR42X1TF U369 ( .A(n485), .B(n498), .C(n1158), .D(n494), .ICI(n1190), .S(
        n482), .ICO(n480), .CO(n481) );
  CMPR42X1TF U370 ( .A(n488), .B(n501), .C(n1094), .D(n497), .ICI(n1126), .S(
        n485), .ICO(n483), .CO(n484) );
  CMPR42X1TF U371 ( .A(n491), .B(n504), .C(n1030), .D(n500), .ICI(n1062), .S(
        n488), .ICO(n486), .CO(n487) );
  CMPR42X1TF U372 ( .A(n493), .B(n506), .C(n966), .D(n503), .ICI(n998), .S(
        n491), .ICO(n489), .CO(n490) );
  CMPR32X2TF U373 ( .A(n1222), .B(n1257), .C(n934), .CO(n492), .S(n493) );
  CMPR42X1TF U374 ( .A(n1159), .B(n499), .C(n508), .D(n1191), .ICI(n1223), .S(
        n496), .ICO(n494), .CO(n495) );
  CMPR42X1TF U375 ( .A(n1095), .B(n502), .C(n511), .D(n1127), .ICI(n512), .S(
        n499), .ICO(n497), .CO(n498) );
  CMPR42X1TF U376 ( .A(n1031), .B(n505), .C(n514), .D(n1063), .ICI(n515), .S(
        n502), .ICO(n500), .CO(n501) );
  CMPR42X1TF U377 ( .A(n967), .B(n507), .C(n517), .D(n999), .ICI(n518), .S(
        n505), .ICO(n503), .CO(n504) );
  CMPR32X2TF U378 ( .A(n935), .B(n7), .C(n520), .CO(n506), .S(n507) );
  CMPR42X1TF U379 ( .A(n1160), .B(n513), .C(n522), .D(n1192), .ICI(n523), .S(
        n510), .ICO(n508), .CO(n509) );
  CMPR42X1TF U380 ( .A(n1096), .B(n516), .C(n525), .D(n1128), .ICI(n526), .S(
        n513), .ICO(n511), .CO(n512) );
  CMPR42X1TF U381 ( .A(n1032), .B(n519), .C(n528), .D(n1064), .ICI(n529), .S(
        n516), .ICO(n514), .CO(n515) );
  CMPR42X1TF U382 ( .A(n968), .B(n521), .C(n531), .D(n1000), .ICI(n532), .S(
        n519), .ICO(n517), .CO(n518) );
  CMPR32X2TF U383 ( .A(n936), .B(n7), .C(n534), .CO(n520), .S(n521) );
  CMPR42X1TF U384 ( .A(n540), .B(n527), .C(n1193), .D(n536), .ICI(n1225), .S(
        n524), .ICO(n522), .CO(n523) );
  CMPR42X1TF U385 ( .A(n543), .B(n530), .C(n1129), .D(n539), .ICI(n1161), .S(
        n527), .ICO(n525), .CO(n526) );
  CMPR42X1TF U386 ( .A(n546), .B(n533), .C(n1065), .D(n542), .ICI(n1097), .S(
        n530), .ICO(n528), .CO(n529) );
  CMPR42X1TF U387 ( .A(n548), .B(n535), .C(n1001), .D(n545), .ICI(n1033), .S(
        n533), .ICO(n531), .CO(n532) );
  CMPR32X2TF U388 ( .A(n937), .B(n7), .C(n969), .CO(n534), .S(n535) );
  CMPR42X1TF U389 ( .A(n541), .B(n1194), .C(n550), .D(n1226), .ICI(n551), .S(
        n538), .ICO(n536), .CO(n537) );
  CMPR42X1TF U390 ( .A(n544), .B(n1130), .C(n553), .D(n1162), .ICI(n554), .S(
        n541), .ICO(n539), .CO(n540) );
  CMPR42X1TF U391 ( .A(n547), .B(n1066), .C(n556), .D(n1098), .ICI(n557), .S(
        n544), .ICO(n542), .CO(n543) );
  CMPR42X1TF U392 ( .A(n549), .B(n1002), .C(n559), .D(n1034), .ICI(n560), .S(
        n547), .ICO(n545), .CO(n546) );
  CMPR32X2TF U393 ( .A(n970), .B(n938), .C(n562), .CO(n548), .S(n549) );
  CMPR42X1TF U394 ( .A(n555), .B(n1195), .C(n564), .D(n1227), .ICI(n565), .S(
        n552), .ICO(n550), .CO(n551) );
  CMPR42X1TF U395 ( .A(n558), .B(n1131), .C(n567), .D(n1163), .ICI(n568), .S(
        n555), .ICO(n553), .CO(n554) );
  CMPR42X1TF U396 ( .A(n561), .B(n1067), .C(n570), .D(n1099), .ICI(n571), .S(
        n558), .ICO(n556), .CO(n557) );
  CMPR42X1TF U397 ( .A(n563), .B(n1003), .C(n573), .D(n1035), .ICI(n574), .S(
        n561), .ICO(n559), .CO(n560) );
  CMPR32X2TF U398 ( .A(n971), .B(n939), .C(n576), .CO(n562), .S(n563) );
  CMPR42X1TF U399 ( .A(n569), .B(n1196), .C(n578), .D(n1228), .ICI(n579), .S(
        n566), .ICO(n564), .CO(n565) );
  CMPR42X1TF U400 ( .A(n572), .B(n1132), .C(n581), .D(n1164), .ICI(n582), .S(
        n569), .ICO(n567), .CO(n568) );
  CMPR42X1TF U401 ( .A(n575), .B(n1068), .C(n584), .D(n1100), .ICI(n585), .S(
        n572), .ICO(n570), .CO(n571) );
  CMPR42X1TF U402 ( .A(n577), .B(n1004), .C(n587), .D(n1036), .ICI(n588), .S(
        n575), .ICO(n573), .CO(n574) );
  CMPR32X2TF U403 ( .A(n972), .B(n940), .C(n590), .CO(n576), .S(n577) );
  CMPR42X1TF U404 ( .A(n583), .B(n1197), .C(n592), .D(n1229), .ICI(n593), .S(
        n580), .ICO(n578), .CO(n579) );
  CMPR42X1TF U405 ( .A(n586), .B(n1133), .C(n595), .D(n1165), .ICI(n596), .S(
        n583), .ICO(n581), .CO(n582) );
  CMPR42X1TF U406 ( .A(n589), .B(n1069), .C(n598), .D(n1101), .ICI(n599), .S(
        n586), .ICO(n584), .CO(n585) );
  CMPR42X1TF U407 ( .A(n591), .B(n1005), .C(n601), .D(n1037), .ICI(n602), .S(
        n589), .ICO(n587), .CO(n588) );
  CMPR32X2TF U408 ( .A(n973), .B(n941), .C(n604), .CO(n590), .S(n591) );
  CMPR42X1TF U409 ( .A(n597), .B(n1198), .C(n606), .D(n1230), .ICI(n607), .S(
        n594), .ICO(n592), .CO(n593) );
  CMPR42X1TF U410 ( .A(n600), .B(n1134), .C(n609), .D(n1166), .ICI(n610), .S(
        n597), .ICO(n595), .CO(n596) );
  CMPR42X1TF U411 ( .A(n603), .B(n1070), .C(n612), .D(n1102), .ICI(n613), .S(
        n600), .ICO(n598), .CO(n599) );
  CMPR42X1TF U412 ( .A(n605), .B(n1006), .C(n615), .D(n1038), .ICI(n616), .S(
        n603), .ICO(n601), .CO(n602) );
  ADDHXLTF U413 ( .A(n974), .B(n618), .CO(n604), .S(n605) );
  CMPR42X1TF U414 ( .A(n611), .B(n1199), .C(n620), .D(n1231), .ICI(n621), .S(
        n608), .ICO(n606), .CO(n607) );
  CMPR42X1TF U415 ( .A(n614), .B(n1135), .C(n623), .D(n1167), .ICI(n624), .S(
        n611), .ICO(n609), .CO(n610) );
  CMPR42X1TF U416 ( .A(n617), .B(n1071), .C(n626), .D(n1103), .ICI(n627), .S(
        n614), .ICO(n612), .CO(n613) );
  CMPR42X1TF U417 ( .A(n619), .B(n1007), .C(n629), .D(n1039), .ICI(n630), .S(
        n617), .ICO(n615), .CO(n616) );
  ADDHXLTF U418 ( .A(n975), .B(n632), .CO(n618), .S(n619) );
  CMPR42X1TF U419 ( .A(n625), .B(n1200), .C(n634), .D(n1232), .ICI(n635), .S(
        n622), .ICO(n620), .CO(n621) );
  CMPR42X1TF U420 ( .A(n628), .B(n1136), .C(n637), .D(n1168), .ICI(n638), .S(
        n625), .ICO(n623), .CO(n624) );
  CMPR42X1TF U421 ( .A(n631), .B(n1072), .C(n640), .D(n1104), .ICI(n641), .S(
        n628), .ICO(n626), .CO(n627) );
  CMPR42X1TF U422 ( .A(n633), .B(n1008), .C(n645), .D(n1040), .ICI(n643), .S(
        n631), .ICO(n629), .CO(n630) );
  ADDHXLTF U423 ( .A(n115), .B(n976), .CO(n632), .S(n633) );
  CMPR42X1TF U424 ( .A(n639), .B(n1201), .C(n647), .D(n1233), .ICI(n648), .S(
        n636), .ICO(n634), .CO(n635) );
  CMPR42X1TF U425 ( .A(n642), .B(n1137), .C(n650), .D(n1169), .ICI(n651), .S(
        n639), .ICO(n637), .CO(n638) );
  CMPR42X1TF U426 ( .A(n644), .B(n1073), .C(n653), .D(n1105), .ICI(n654), .S(
        n642), .ICO(n640), .CO(n641) );
  CMPR32X2TF U427 ( .A(n1041), .B(n646), .C(n656), .CO(n643), .S(n644) );
  ADDHXLTF U428 ( .A(n1009), .B(n658), .CO(n645), .S(n646) );
  CMPR42X1TF U429 ( .A(n652), .B(n1202), .C(n660), .D(n1234), .ICI(n661), .S(
        n649), .ICO(n647), .CO(n648) );
  CMPR42X1TF U430 ( .A(n655), .B(n1138), .C(n663), .D(n1170), .ICI(n664), .S(
        n652), .ICO(n650), .CO(n651) );
  CMPR42X1TF U431 ( .A(n657), .B(n1074), .C(n666), .D(n1106), .ICI(n667), .S(
        n655), .ICO(n653), .CO(n654) );
  CMPR32X2TF U432 ( .A(n1042), .B(n659), .C(n669), .CO(n656), .S(n657) );
  ADDHXLTF U433 ( .A(n1010), .B(n671), .CO(n658), .S(n659) );
  CMPR42X1TF U434 ( .A(n665), .B(n1203), .C(n673), .D(n1235), .ICI(n674), .S(
        n662), .ICO(n660), .CO(n661) );
  CMPR42X1TF U435 ( .A(n668), .B(n1139), .C(n676), .D(n1171), .ICI(n677), .S(
        n665), .ICO(n663), .CO(n664) );
  CMPR42X1TF U436 ( .A(n670), .B(n1075), .C(n679), .D(n1107), .ICI(n680), .S(
        n668), .ICO(n666), .CO(n667) );
  CMPR32X2TF U437 ( .A(n1043), .B(n672), .C(n682), .CO(n669), .S(n670) );
  ADDHXLTF U438 ( .A(n103), .B(n1011), .CO(n671), .S(n672) );
  CMPR42X1TF U439 ( .A(n678), .B(n1204), .C(n684), .D(n1236), .ICI(n685), .S(
        n675), .ICO(n673), .CO(n674) );
  CMPR42X1TF U440 ( .A(n681), .B(n1140), .C(n687), .D(n1172), .ICI(n688), .S(
        n678), .ICO(n676), .CO(n677) );
  CMPR42X1TF U441 ( .A(n683), .B(n1076), .C(n690), .D(n1108), .ICI(n691), .S(
        n681), .ICO(n679), .CO(n680) );
  ADDHXLTF U442 ( .A(n1044), .B(n693), .CO(n682), .S(n683) );
  CMPR42X1TF U443 ( .A(n689), .B(n1205), .C(n695), .D(n1237), .ICI(n696), .S(
        n686), .ICO(n684), .CO(n685) );
  CMPR42X1TF U444 ( .A(n692), .B(n1141), .C(n698), .D(n1173), .ICI(n699), .S(
        n689), .ICO(n687), .CO(n688) );
  CMPR42X1TF U445 ( .A(n694), .B(n1077), .C(n701), .D(n1109), .ICI(n702), .S(
        n692), .ICO(n690), .CO(n691) );
  ADDHXLTF U446 ( .A(n1045), .B(n704), .CO(n693), .S(n694) );
  CMPR42X1TF U447 ( .A(n700), .B(n1206), .C(n706), .D(n1238), .ICI(n707), .S(
        n697), .ICO(n695), .CO(n696) );
  CMPR42X1TF U448 ( .A(n703), .B(n1142), .C(n709), .D(n1174), .ICI(n710), .S(
        n700), .ICO(n698), .CO(n699) );
  CMPR42X1TF U449 ( .A(n705), .B(n1078), .C(n714), .D(n1110), .ICI(n712), .S(
        n703), .ICO(n701), .CO(n702) );
  ADDHXLTF U450 ( .A(n91), .B(n1046), .CO(n704), .S(n705) );
  CMPR42X1TF U451 ( .A(n711), .B(n1207), .C(n716), .D(n1239), .ICI(n717), .S(
        n708), .ICO(n706), .CO(n707) );
  CMPR42X1TF U452 ( .A(n713), .B(n1143), .C(n719), .D(n1175), .ICI(n720), .S(
        n711), .ICO(n709), .CO(n710) );
  CMPR32X2TF U453 ( .A(n1111), .B(n715), .C(n722), .CO(n712), .S(n713) );
  ADDHXLTF U454 ( .A(n1079), .B(n724), .CO(n714), .S(n715) );
  CMPR42X1TF U455 ( .A(n721), .B(n1208), .C(n726), .D(n1240), .ICI(n727), .S(
        n718), .ICO(n716), .CO(n717) );
  CMPR42X1TF U456 ( .A(n723), .B(n1144), .C(n729), .D(n1176), .ICI(n730), .S(
        n721), .ICO(n719), .CO(n720) );
  CMPR32X2TF U457 ( .A(n1112), .B(n725), .C(n732), .CO(n722), .S(n723) );
  ADDHXLTF U458 ( .A(n1080), .B(n734), .CO(n724), .S(n725) );
  CMPR42X1TF U459 ( .A(n731), .B(n1209), .C(n736), .D(n1241), .ICI(n737), .S(
        n728), .ICO(n726), .CO(n727) );
  CMPR42X1TF U460 ( .A(n733), .B(n1145), .C(n739), .D(n1177), .ICI(n740), .S(
        n731), .ICO(n729), .CO(n730) );
  CMPR32X2TF U461 ( .A(n1113), .B(n735), .C(n742), .CO(n732), .S(n733) );
  ADDHXLTF U462 ( .A(n79), .B(n1081), .CO(n734), .S(n735) );
  CMPR42X1TF U463 ( .A(n741), .B(n1210), .C(n744), .D(n1242), .ICI(n745), .S(
        n738), .ICO(n736), .CO(n737) );
  CMPR42X1TF U464 ( .A(n743), .B(n1146), .C(n747), .D(n1178), .ICI(n748), .S(
        n741), .ICO(n739), .CO(n740) );
  ADDHXLTF U465 ( .A(n1114), .B(n750), .CO(n742), .S(n743) );
  CMPR42X1TF U466 ( .A(n749), .B(n1211), .C(n752), .D(n1243), .ICI(n753), .S(
        n746), .ICO(n744), .CO(n745) );
  CMPR42X1TF U467 ( .A(n751), .B(n1147), .C(n755), .D(n1179), .ICI(n756), .S(
        n749), .ICO(n747), .CO(n748) );
  ADDHXLTF U468 ( .A(n1115), .B(n758), .CO(n750), .S(n751) );
  CMPR42X1TF U469 ( .A(n757), .B(n1212), .C(n760), .D(n1244), .ICI(n761), .S(
        n754), .ICO(n752), .CO(n753) );
  CMPR42X1TF U470 ( .A(n759), .B(n1148), .C(n765), .D(n1180), .ICI(n763), .S(
        n757), .ICO(n755), .CO(n756) );
  ADDHXLTF U471 ( .A(n67), .B(n1116), .CO(n758), .S(n759) );
  CMPR42X1TF U472 ( .A(n764), .B(n1213), .C(n767), .D(n1245), .ICI(n768), .S(
        n762), .ICO(n760), .CO(n761) );
  CMPR32X2TF U473 ( .A(n1181), .B(n766), .C(n770), .CO(n763), .S(n764) );
  ADDHXLTF U474 ( .A(n1149), .B(n772), .CO(n765), .S(n766) );
  CMPR42X1TF U475 ( .A(n771), .B(n1214), .C(n774), .D(n1246), .ICI(n775), .S(
        n769), .ICO(n767), .CO(n768) );
  CMPR32X2TF U476 ( .A(n1182), .B(n773), .C(n777), .CO(n770), .S(n771) );
  ADDHXLTF U477 ( .A(n1150), .B(n779), .CO(n772), .S(n773) );
  CMPR42X1TF U478 ( .A(n778), .B(n1215), .C(n781), .D(n1247), .ICI(n782), .S(
        n776), .ICO(n774), .CO(n775) );
  CMPR32X2TF U479 ( .A(n1183), .B(n780), .C(n784), .CO(n777), .S(n778) );
  ADDHXLTF U480 ( .A(n55), .B(n1151), .CO(n779), .S(n780) );
  CMPR42X1TF U481 ( .A(n785), .B(n1216), .C(n786), .D(n1248), .ICI(n787), .S(
        n783), .ICO(n781), .CO(n782) );
  ADDHXLTF U482 ( .A(n1184), .B(n789), .CO(n784), .S(n785) );
  CMPR42X1TF U483 ( .A(n790), .B(n1217), .C(n791), .D(n1249), .ICI(n792), .S(
        n788), .ICO(n786), .CO(n787) );
  ADDHXLTF U484 ( .A(n1185), .B(n794), .CO(n789), .S(n790) );
  CMPR42X1TF U485 ( .A(n795), .B(n1218), .C(n798), .D(n1250), .ICI(n796), .S(
        n793), .ICO(n791), .CO(n792) );
  ADDHXLTF U486 ( .A(n43), .B(n1186), .CO(n794), .S(n795) );
  CMPR32X2TF U487 ( .A(n1251), .B(n799), .C(n800), .CO(n796), .S(n797) );
  ADDHXLTF U488 ( .A(n1219), .B(n802), .CO(n798), .S(n799) );
  CMPR32X2TF U489 ( .A(n1252), .B(n803), .C(n804), .CO(n800), .S(n801) );
  ADDHXLTF U490 ( .A(n1220), .B(n806), .CO(n802), .S(n803) );
  CMPR32X2TF U491 ( .A(n1253), .B(n807), .C(n808), .CO(n804), .S(n805) );
  ADDHXLTF U492 ( .A(n31), .B(n1221), .CO(n806), .S(n807) );
  ADDHXLTF U493 ( .A(n1254), .B(n810), .CO(n808), .S(n809) );
  ADDHXLTF U494 ( .A(n1255), .B(n812), .CO(n810), .S(n811) );
  ADDHXLTF U495 ( .A(n19), .B(n1256), .CO(n812), .S(n813) );
  NAND2X1TF U497 ( .A(n129), .B(n225), .Y(n1292) );
  OAI21X1TF U498 ( .A0(n2007), .A1(n127), .B0(n1293), .Y(n291) );
  AOI21X1TF U499 ( .A0(n129), .A1(n222), .B0(n814), .Y(n1293) );
  AND2X2TF U500 ( .A(n124), .B(n225), .Y(n814) );
  OAI21X1TF U501 ( .A0(n2008), .A1(n127), .B0(n1294), .Y(n913) );
  AOI222XLTF U502 ( .A0(n122), .A1(n225), .B0(n124), .B1(n222), .C0(n129), 
        .C1(n219), .Y(n1294) );
  OAI21X1TF U503 ( .A0(n2009), .A1(n127), .B0(n1295), .Y(n914) );
  AOI222XLTF U504 ( .A0(n122), .A1(n222), .B0(n124), .B1(n219), .C0(n129), 
        .C1(n216), .Y(n1295) );
  OAI21X1TF U505 ( .A0(n2010), .A1(n127), .B0(n1296), .Y(n915) );
  AOI222XLTF U506 ( .A0(n122), .A1(n219), .B0(n124), .B1(n216), .C0(n129), 
        .C1(n213), .Y(n1296) );
  OAI21X1TF U507 ( .A0(n2011), .A1(n127), .B0(n1297), .Y(n916) );
  AOI222XLTF U508 ( .A0(n122), .A1(n216), .B0(n124), .B1(n213), .C0(n129), 
        .C1(n210), .Y(n1297) );
  OAI21X1TF U509 ( .A0(n2012), .A1(n127), .B0(n1298), .Y(n917) );
  AOI222XLTF U510 ( .A0(n122), .A1(n213), .B0(n124), .B1(n210), .C0(n129), 
        .C1(n207), .Y(n1298) );
  OAI21X1TF U511 ( .A0(n2013), .A1(n127), .B0(n1299), .Y(n918) );
  AOI222XLTF U512 ( .A0(n122), .A1(n210), .B0(n124), .B1(n207), .C0(n129), 
        .C1(n204), .Y(n1299) );
  OAI21X1TF U513 ( .A0(n2014), .A1(n127), .B0(n1300), .Y(n919) );
  AOI222XLTF U514 ( .A0(n122), .A1(n207), .B0(n124), .B1(n204), .C0(n129), 
        .C1(n201), .Y(n1300) );
  OAI21X1TF U515 ( .A0(n2015), .A1(n127), .B0(n1301), .Y(n920) );
  AOI222XLTF U516 ( .A0(n122), .A1(n204), .B0(n124), .B1(n201), .C0(n129), 
        .C1(n198), .Y(n1301) );
  OAI21X1TF U517 ( .A0(n2016), .A1(n127), .B0(n1302), .Y(n921) );
  AOI222XLTF U518 ( .A0(n122), .A1(n201), .B0(n124), .B1(n198), .C0(n129), 
        .C1(n195), .Y(n1302) );
  OAI21X1TF U519 ( .A0(n2017), .A1(n127), .B0(n1303), .Y(n922) );
  AOI222XLTF U520 ( .A0(n122), .A1(n198), .B0(n124), .B1(n195), .C0(n129), 
        .C1(n192), .Y(n1303) );
  OAI21X1TF U521 ( .A0(n2018), .A1(n126), .B0(n1304), .Y(n923) );
  AOI222XLTF U522 ( .A0(n122), .A1(n195), .B0(n124), .B1(n192), .C0(n129), 
        .C1(n189), .Y(n1304) );
  OAI21X1TF U523 ( .A0(n2019), .A1(n126), .B0(n1305), .Y(n341) );
  AOI222XLTF U524 ( .A0(n122), .A1(n192), .B0(n124), .B1(n189), .C0(n129), 
        .C1(n186), .Y(n1305) );
  OAI21X1TF U525 ( .A0(n2020), .A1(n126), .B0(n1306), .Y(n924) );
  AOI222XLTF U526 ( .A0(n122), .A1(n189), .B0(n124), .B1(n186), .C0(n129), 
        .C1(n183), .Y(n1306) );
  OAI21X1TF U527 ( .A0(n2021), .A1(n126), .B0(n1307), .Y(n925) );
  AOI222XLTF U528 ( .A0(n122), .A1(n186), .B0(n124), .B1(n183), .C0(n129), 
        .C1(n180), .Y(n1307) );
  OAI21X1TF U529 ( .A0(n2022), .A1(n126), .B0(n1308), .Y(n926) );
  AOI222XLTF U530 ( .A0(n122), .A1(n183), .B0(n124), .B1(n180), .C0(n128), 
        .C1(n177), .Y(n1308) );
  OAI21X1TF U531 ( .A0(n2023), .A1(n126), .B0(n1309), .Y(n927) );
  AOI222XLTF U532 ( .A0(n122), .A1(n180), .B0(n123), .B1(n177), .C0(n128), 
        .C1(n174), .Y(n1309) );
  OAI21X1TF U533 ( .A0(n2024), .A1(n126), .B0(n1310), .Y(n928) );
  AOI222XLTF U534 ( .A0(n121), .A1(n177), .B0(n123), .B1(n174), .C0(n128), 
        .C1(n171), .Y(n1310) );
  OAI21X1TF U535 ( .A0(n2025), .A1(n126), .B0(n1311), .Y(n394) );
  AOI222XLTF U536 ( .A0(n121), .A1(n174), .B0(n123), .B1(n171), .C0(n128), 
        .C1(n168), .Y(n1311) );
  OAI21X1TF U537 ( .A0(n2026), .A1(n126), .B0(n1312), .Y(n929) );
  AOI222XLTF U538 ( .A0(n121), .A1(n171), .B0(n123), .B1(n168), .C0(n128), 
        .C1(n165), .Y(n1312) );
  OAI21X1TF U539 ( .A0(n2027), .A1(n126), .B0(n1313), .Y(n930) );
  AOI222XLTF U540 ( .A0(n121), .A1(n168), .B0(n123), .B1(n165), .C0(n128), 
        .C1(n162), .Y(n1313) );
  OAI21X1TF U541 ( .A0(n2028), .A1(n126), .B0(n1314), .Y(n931) );
  AOI222XLTF U542 ( .A0(n121), .A1(n165), .B0(n123), .B1(n162), .C0(n128), 
        .C1(n159), .Y(n1314) );
  OAI21X1TF U543 ( .A0(n2029), .A1(n126), .B0(n1315), .Y(n932) );
  AOI222XLTF U544 ( .A0(n121), .A1(n162), .B0(n123), .B1(n159), .C0(n128), 
        .C1(n156), .Y(n1315) );
  OAI21X1TF U545 ( .A0(n2030), .A1(n125), .B0(n1316), .Y(n933) );
  AOI222XLTF U546 ( .A0(n121), .A1(n159), .B0(n123), .B1(n156), .C0(n128), 
        .C1(n153), .Y(n1316) );
  OAI21X1TF U547 ( .A0(n2031), .A1(n125), .B0(n1317), .Y(n465) );
  AOI222XLTF U548 ( .A0(n121), .A1(n156), .B0(n123), .B1(n153), .C0(n128), 
        .C1(n150), .Y(n1317) );
  OAI21X1TF U549 ( .A0(n2032), .A1(n125), .B0(n1318), .Y(n934) );
  AOI222XLTF U550 ( .A0(n121), .A1(n153), .B0(n123), .B1(n150), .C0(n128), 
        .C1(n147), .Y(n1318) );
  OAI21X1TF U551 ( .A0(n2033), .A1(n125), .B0(n1319), .Y(n935) );
  AOI222XLTF U552 ( .A0(n121), .A1(n150), .B0(n123), .B1(n147), .C0(n128), 
        .C1(n144), .Y(n1319) );
  OAI21X1TF U553 ( .A0(n2034), .A1(n125), .B0(n1320), .Y(n936) );
  AOI222XLTF U554 ( .A0(n121), .A1(n147), .B0(n123), .B1(n144), .C0(n128), 
        .C1(n141), .Y(n1320) );
  OAI21X1TF U555 ( .A0(n2035), .A1(n125), .B0(n1321), .Y(n937) );
  AOI222XLTF U556 ( .A0(n121), .A1(n144), .B0(n123), .B1(n141), .C0(n128), 
        .C1(n138), .Y(n1321) );
  OAI21X1TF U557 ( .A0(n2036), .A1(n125), .B0(n1322), .Y(n938) );
  AOI222XLTF U558 ( .A0(n121), .A1(n141), .B0(n123), .B1(n138), .C0(n128), 
        .C1(n135), .Y(n1322) );
  OAI21X1TF U559 ( .A0(n2037), .A1(n125), .B0(n1323), .Y(n939) );
  AOI222XLTF U560 ( .A0(n121), .A1(n138), .B0(n123), .B1(n135), .C0(n128), 
        .C1(n132), .Y(n1323) );
  OAI21X1TF U561 ( .A0(n125), .A1(n2038), .B0(n2300), .Y(n940) );
  OAI21X1TF U564 ( .A0(n125), .A1(n2039), .B0(n2311), .Y(n941) );
  INVX2TF U567 ( .A(n115), .Y(n942) );
  XOR2X1TF U568 ( .A(n1326), .B(n115), .Y(n943) );
  OAI21X1TF U569 ( .A0(n2006), .A1(n118), .B0(n1360), .Y(n1326) );
  NAND2X1TF U570 ( .A(n120), .B(n225), .Y(n1360) );
  XOR2X1TF U571 ( .A(n1327), .B(n115), .Y(n944) );
  OAI21X1TF U572 ( .A0(n2007), .A1(n118), .B0(n1361), .Y(n1327) );
  AOI21X1TF U573 ( .A0(n120), .A1(n222), .B0(n817), .Y(n1361) );
  AND2X2TF U574 ( .A(n112), .B(n225), .Y(n817) );
  XOR2X1TF U575 ( .A(n1328), .B(n115), .Y(n945) );
  OAI21X1TF U576 ( .A0(n2008), .A1(n118), .B0(n1362), .Y(n1328) );
  AOI222XLTF U577 ( .A0(n110), .A1(n225), .B0(n112), .B1(n222), .C0(n120), 
        .C1(n219), .Y(n1362) );
  XOR2X1TF U578 ( .A(n1329), .B(n115), .Y(n946) );
  OAI21X1TF U579 ( .A0(n2009), .A1(n118), .B0(n1363), .Y(n1329) );
  AOI222XLTF U580 ( .A0(n110), .A1(n222), .B0(n112), .B1(n219), .C0(n120), 
        .C1(n216), .Y(n1363) );
  XOR2X1TF U581 ( .A(n1330), .B(n115), .Y(n947) );
  OAI21X1TF U582 ( .A0(n2010), .A1(n118), .B0(n1364), .Y(n1330) );
  AOI222XLTF U583 ( .A0(n110), .A1(n219), .B0(n112), .B1(n216), .C0(n120), 
        .C1(n213), .Y(n1364) );
  XOR2X1TF U584 ( .A(n1331), .B(n115), .Y(n948) );
  OAI21X1TF U585 ( .A0(n2011), .A1(n118), .B0(n1365), .Y(n1331) );
  AOI222XLTF U586 ( .A0(n110), .A1(n216), .B0(n112), .B1(n213), .C0(n120), 
        .C1(n210), .Y(n1365) );
  XOR2X1TF U587 ( .A(n1332), .B(n115), .Y(n949) );
  OAI21X1TF U588 ( .A0(n2012), .A1(n118), .B0(n1366), .Y(n1332) );
  AOI222XLTF U589 ( .A0(n110), .A1(n213), .B0(n112), .B1(n210), .C0(n120), 
        .C1(n207), .Y(n1366) );
  XOR2X1TF U590 ( .A(n1333), .B(n115), .Y(n950) );
  OAI21X1TF U591 ( .A0(n2013), .A1(n118), .B0(n1367), .Y(n1333) );
  AOI222XLTF U592 ( .A0(n110), .A1(n210), .B0(n112), .B1(n207), .C0(n120), 
        .C1(n204), .Y(n1367) );
  XOR2X1TF U593 ( .A(n1334), .B(n115), .Y(n951) );
  OAI21X1TF U594 ( .A0(n2014), .A1(n118), .B0(n1368), .Y(n1334) );
  AOI222XLTF U595 ( .A0(n110), .A1(n207), .B0(n112), .B1(n204), .C0(n120), 
        .C1(n201), .Y(n1368) );
  XOR2X1TF U596 ( .A(n1335), .B(n115), .Y(n952) );
  OAI21X1TF U597 ( .A0(n2015), .A1(n118), .B0(n1369), .Y(n1335) );
  AOI222XLTF U598 ( .A0(n110), .A1(n204), .B0(n112), .B1(n201), .C0(n120), 
        .C1(n198), .Y(n1369) );
  XOR2X1TF U599 ( .A(n1336), .B(n114), .Y(n953) );
  OAI21X1TF U600 ( .A0(n2016), .A1(n118), .B0(n1370), .Y(n1336) );
  AOI222XLTF U601 ( .A0(n110), .A1(n201), .B0(n112), .B1(n198), .C0(n120), 
        .C1(n195), .Y(n1370) );
  XOR2X1TF U602 ( .A(n1337), .B(n114), .Y(n954) );
  OAI21X1TF U603 ( .A0(n2017), .A1(n118), .B0(n1371), .Y(n1337) );
  AOI222XLTF U604 ( .A0(n110), .A1(n198), .B0(n112), .B1(n195), .C0(n120), 
        .C1(n192), .Y(n1371) );
  XOR2X1TF U605 ( .A(n1338), .B(n114), .Y(n955) );
  OAI21X1TF U606 ( .A0(n2018), .A1(n117), .B0(n1372), .Y(n1338) );
  AOI222XLTF U607 ( .A0(n110), .A1(n195), .B0(n112), .B1(n192), .C0(n120), 
        .C1(n189), .Y(n1372) );
  XOR2X1TF U608 ( .A(n1339), .B(n114), .Y(n956) );
  OAI21X1TF U609 ( .A0(n2019), .A1(n117), .B0(n1373), .Y(n1339) );
  AOI222XLTF U610 ( .A0(n110), .A1(n192), .B0(n112), .B1(n189), .C0(n120), 
        .C1(n186), .Y(n1373) );
  XOR2X1TF U611 ( .A(n1340), .B(n114), .Y(n957) );
  OAI21X1TF U612 ( .A0(n2020), .A1(n117), .B0(n1374), .Y(n1340) );
  AOI222XLTF U613 ( .A0(n110), .A1(n189), .B0(n112), .B1(n186), .C0(n120), 
        .C1(n183), .Y(n1374) );
  XOR2X1TF U614 ( .A(n1341), .B(n114), .Y(n958) );
  OAI21X1TF U615 ( .A0(n2021), .A1(n117), .B0(n1375), .Y(n1341) );
  AOI222XLTF U616 ( .A0(n110), .A1(n186), .B0(n112), .B1(n183), .C0(n120), 
        .C1(n180), .Y(n1375) );
  XOR2X1TF U617 ( .A(n1342), .B(n114), .Y(n959) );
  OAI21X1TF U618 ( .A0(n2022), .A1(n117), .B0(n1376), .Y(n1342) );
  AOI222XLTF U619 ( .A0(n110), .A1(n183), .B0(n112), .B1(n180), .C0(n119), 
        .C1(n177), .Y(n1376) );
  XOR2X1TF U620 ( .A(n1343), .B(n114), .Y(n960) );
  OAI21X1TF U621 ( .A0(n2023), .A1(n117), .B0(n1377), .Y(n1343) );
  AOI222XLTF U622 ( .A0(n110), .A1(n180), .B0(n111), .B1(n177), .C0(n119), 
        .C1(n174), .Y(n1377) );
  XOR2X1TF U623 ( .A(n1344), .B(n114), .Y(n961) );
  OAI21X1TF U624 ( .A0(n2024), .A1(n117), .B0(n1378), .Y(n1344) );
  AOI222XLTF U625 ( .A0(n109), .A1(n177), .B0(n111), .B1(n174), .C0(n119), 
        .C1(n171), .Y(n1378) );
  XOR2X1TF U626 ( .A(n1345), .B(n114), .Y(n962) );
  OAI21X1TF U627 ( .A0(n2025), .A1(n117), .B0(n1379), .Y(n1345) );
  AOI222XLTF U628 ( .A0(n109), .A1(n174), .B0(n111), .B1(n171), .C0(n119), 
        .C1(n168), .Y(n1379) );
  XOR2X1TF U629 ( .A(n1346), .B(n114), .Y(n963) );
  OAI21X1TF U630 ( .A0(n2026), .A1(n117), .B0(n1380), .Y(n1346) );
  AOI222XLTF U631 ( .A0(n109), .A1(n171), .B0(n111), .B1(n168), .C0(n119), 
        .C1(n165), .Y(n1380) );
  XOR2X1TF U632 ( .A(n1347), .B(n114), .Y(n964) );
  OAI21X1TF U633 ( .A0(n2027), .A1(n117), .B0(n1381), .Y(n1347) );
  AOI222XLTF U634 ( .A0(n109), .A1(n168), .B0(n111), .B1(n165), .C0(n119), 
        .C1(n162), .Y(n1381) );
  XOR2X1TF U635 ( .A(n1348), .B(n113), .Y(n965) );
  OAI21X1TF U636 ( .A0(n2028), .A1(n117), .B0(n1382), .Y(n1348) );
  AOI222XLTF U637 ( .A0(n109), .A1(n165), .B0(n111), .B1(n162), .C0(n119), 
        .C1(n159), .Y(n1382) );
  XOR2X1TF U638 ( .A(n1349), .B(n113), .Y(n966) );
  OAI21X1TF U639 ( .A0(n2029), .A1(n117), .B0(n1383), .Y(n1349) );
  AOI222XLTF U640 ( .A0(n109), .A1(n162), .B0(n111), .B1(n159), .C0(n119), 
        .C1(n156), .Y(n1383) );
  XOR2X1TF U641 ( .A(n1350), .B(n113), .Y(n967) );
  OAI21X1TF U642 ( .A0(n2030), .A1(n116), .B0(n1384), .Y(n1350) );
  AOI222XLTF U643 ( .A0(n109), .A1(n159), .B0(n111), .B1(n156), .C0(n119), 
        .C1(n153), .Y(n1384) );
  XOR2X1TF U644 ( .A(n1351), .B(n113), .Y(n968) );
  OAI21X1TF U645 ( .A0(n2031), .A1(n116), .B0(n1385), .Y(n1351) );
  AOI222XLTF U646 ( .A0(n109), .A1(n156), .B0(n111), .B1(n153), .C0(n119), 
        .C1(n150), .Y(n1385) );
  XOR2X1TF U647 ( .A(n1352), .B(n113), .Y(n969) );
  OAI21X1TF U648 ( .A0(n2032), .A1(n116), .B0(n1386), .Y(n1352) );
  AOI222XLTF U649 ( .A0(n109), .A1(n153), .B0(n111), .B1(n150), .C0(n119), 
        .C1(n147), .Y(n1386) );
  XOR2X1TF U650 ( .A(n1353), .B(n113), .Y(n970) );
  OAI21X1TF U651 ( .A0(n2033), .A1(n116), .B0(n1387), .Y(n1353) );
  AOI222XLTF U652 ( .A0(n109), .A1(n150), .B0(n111), .B1(n147), .C0(n119), 
        .C1(n144), .Y(n1387) );
  XOR2X1TF U653 ( .A(n1354), .B(n113), .Y(n971) );
  OAI21X1TF U654 ( .A0(n2034), .A1(n116), .B0(n1388), .Y(n1354) );
  AOI222XLTF U655 ( .A0(n109), .A1(n147), .B0(n111), .B1(n144), .C0(n119), 
        .C1(n141), .Y(n1388) );
  XOR2X1TF U656 ( .A(n1355), .B(n113), .Y(n972) );
  OAI21X1TF U657 ( .A0(n2035), .A1(n116), .B0(n1389), .Y(n1355) );
  AOI222XLTF U658 ( .A0(n109), .A1(n144), .B0(n111), .B1(n141), .C0(n119), 
        .C1(n138), .Y(n1389) );
  XOR2X1TF U659 ( .A(n1356), .B(n113), .Y(n973) );
  OAI21X1TF U660 ( .A0(n2036), .A1(n116), .B0(n1390), .Y(n1356) );
  AOI222XLTF U661 ( .A0(n109), .A1(n141), .B0(n111), .B1(n138), .C0(n119), 
        .C1(n135), .Y(n1390) );
  XOR2X1TF U662 ( .A(n1357), .B(n113), .Y(n974) );
  OAI21X1TF U663 ( .A0(n2037), .A1(n116), .B0(n1391), .Y(n1357) );
  AOI222XLTF U664 ( .A0(n109), .A1(n138), .B0(n111), .B1(n135), .C0(n119), 
        .C1(n132), .Y(n1391) );
  XOR2X1TF U665 ( .A(n1358), .B(n113), .Y(n975) );
  OAI21X1TF U666 ( .A0(n116), .A1(n2038), .B0(n2299), .Y(n1358) );
  XOR2X1TF U669 ( .A(n1359), .B(n113), .Y(n976) );
  OAI21X1TF U670 ( .A0(n116), .A1(n2039), .B0(n2310), .Y(n1359) );
  INVX2TF U673 ( .A(n103), .Y(n977) );
  XOR2X1TF U674 ( .A(n1394), .B(n103), .Y(n978) );
  OAI21X1TF U675 ( .A0(n2006), .A1(n106), .B0(n1428), .Y(n1394) );
  NAND2X1TF U676 ( .A(n108), .B(n225), .Y(n1428) );
  XOR2X1TF U677 ( .A(n1395), .B(n103), .Y(n979) );
  OAI21X1TF U678 ( .A0(n2007), .A1(n106), .B0(n1429), .Y(n1395) );
  AOI21X1TF U679 ( .A0(n108), .A1(n222), .B0(n820), .Y(n1429) );
  AND2X2TF U680 ( .A(n100), .B(n225), .Y(n820) );
  XOR2X1TF U681 ( .A(n1396), .B(n103), .Y(n980) );
  OAI21X1TF U682 ( .A0(n2008), .A1(n106), .B0(n1430), .Y(n1396) );
  AOI222XLTF U683 ( .A0(n98), .A1(n225), .B0(n100), .B1(n222), .C0(n108), .C1(
        n219), .Y(n1430) );
  XOR2X1TF U684 ( .A(n1397), .B(n103), .Y(n981) );
  OAI21X1TF U685 ( .A0(n2009), .A1(n106), .B0(n1431), .Y(n1397) );
  AOI222XLTF U686 ( .A0(n98), .A1(n222), .B0(n100), .B1(n219), .C0(n108), .C1(
        n216), .Y(n1431) );
  XOR2X1TF U687 ( .A(n1398), .B(n103), .Y(n982) );
  OAI21X1TF U688 ( .A0(n2010), .A1(n106), .B0(n1432), .Y(n1398) );
  AOI222XLTF U689 ( .A0(n98), .A1(n219), .B0(n100), .B1(n216), .C0(n108), .C1(
        n213), .Y(n1432) );
  XOR2X1TF U690 ( .A(n1399), .B(n103), .Y(n983) );
  OAI21X1TF U691 ( .A0(n2011), .A1(n106), .B0(n1433), .Y(n1399) );
  AOI222XLTF U692 ( .A0(n98), .A1(n216), .B0(n100), .B1(n213), .C0(n108), .C1(
        n210), .Y(n1433) );
  XOR2X1TF U693 ( .A(n1400), .B(n103), .Y(n984) );
  OAI21X1TF U694 ( .A0(n2012), .A1(n106), .B0(n1434), .Y(n1400) );
  AOI222XLTF U695 ( .A0(n98), .A1(n213), .B0(n100), .B1(n210), .C0(n108), .C1(
        n207), .Y(n1434) );
  XOR2X1TF U696 ( .A(n1401), .B(n103), .Y(n985) );
  OAI21X1TF U697 ( .A0(n2013), .A1(n106), .B0(n1435), .Y(n1401) );
  AOI222XLTF U698 ( .A0(n98), .A1(n210), .B0(n100), .B1(n207), .C0(n108), .C1(
        n204), .Y(n1435) );
  XOR2X1TF U699 ( .A(n1402), .B(n103), .Y(n986) );
  OAI21X1TF U700 ( .A0(n2014), .A1(n106), .B0(n1436), .Y(n1402) );
  AOI222XLTF U701 ( .A0(n98), .A1(n207), .B0(n100), .B1(n204), .C0(n108), .C1(
        n201), .Y(n1436) );
  XOR2X1TF U702 ( .A(n1403), .B(n103), .Y(n987) );
  OAI21X1TF U703 ( .A0(n2015), .A1(n106), .B0(n1437), .Y(n1403) );
  AOI222XLTF U704 ( .A0(n98), .A1(n204), .B0(n100), .B1(n201), .C0(n108), .C1(
        n198), .Y(n1437) );
  XOR2X1TF U705 ( .A(n1404), .B(n102), .Y(n988) );
  OAI21X1TF U706 ( .A0(n2016), .A1(n106), .B0(n1438), .Y(n1404) );
  AOI222XLTF U707 ( .A0(n98), .A1(n201), .B0(n100), .B1(n198), .C0(n108), .C1(
        n195), .Y(n1438) );
  XOR2X1TF U708 ( .A(n1405), .B(n102), .Y(n989) );
  OAI21X1TF U709 ( .A0(n2017), .A1(n106), .B0(n1439), .Y(n1405) );
  AOI222XLTF U710 ( .A0(n98), .A1(n198), .B0(n100), .B1(n195), .C0(n108), .C1(
        n192), .Y(n1439) );
  XOR2X1TF U711 ( .A(n1406), .B(n102), .Y(n990) );
  OAI21X1TF U712 ( .A0(n2018), .A1(n105), .B0(n1440), .Y(n1406) );
  AOI222XLTF U713 ( .A0(n98), .A1(n195), .B0(n100), .B1(n192), .C0(n108), .C1(
        n189), .Y(n1440) );
  XOR2X1TF U714 ( .A(n1407), .B(n102), .Y(n991) );
  OAI21X1TF U715 ( .A0(n2019), .A1(n105), .B0(n1441), .Y(n1407) );
  AOI222XLTF U716 ( .A0(n98), .A1(n192), .B0(n100), .B1(n189), .C0(n108), .C1(
        n186), .Y(n1441) );
  XOR2X1TF U717 ( .A(n1408), .B(n102), .Y(n992) );
  OAI21X1TF U718 ( .A0(n2020), .A1(n105), .B0(n1442), .Y(n1408) );
  AOI222XLTF U719 ( .A0(n98), .A1(n189), .B0(n100), .B1(n186), .C0(n108), .C1(
        n183), .Y(n1442) );
  XOR2X1TF U720 ( .A(n1409), .B(n102), .Y(n993) );
  OAI21X1TF U721 ( .A0(n2021), .A1(n105), .B0(n1443), .Y(n1409) );
  AOI222XLTF U722 ( .A0(n98), .A1(n186), .B0(n100), .B1(n183), .C0(n108), .C1(
        n180), .Y(n1443) );
  XOR2X1TF U723 ( .A(n1410), .B(n102), .Y(n994) );
  OAI21X1TF U724 ( .A0(n2022), .A1(n105), .B0(n1444), .Y(n1410) );
  AOI222XLTF U725 ( .A0(n98), .A1(n183), .B0(n100), .B1(n180), .C0(n107), .C1(
        n177), .Y(n1444) );
  XOR2X1TF U726 ( .A(n1411), .B(n102), .Y(n995) );
  OAI21X1TF U727 ( .A0(n2023), .A1(n105), .B0(n1445), .Y(n1411) );
  AOI222XLTF U728 ( .A0(n98), .A1(n180), .B0(n99), .B1(n177), .C0(n107), .C1(
        n174), .Y(n1445) );
  XOR2X1TF U729 ( .A(n1412), .B(n102), .Y(n996) );
  OAI21X1TF U730 ( .A0(n2024), .A1(n105), .B0(n1446), .Y(n1412) );
  AOI222XLTF U731 ( .A0(n97), .A1(n177), .B0(n99), .B1(n174), .C0(n107), .C1(
        n171), .Y(n1446) );
  XOR2X1TF U732 ( .A(n1413), .B(n102), .Y(n997) );
  OAI21X1TF U733 ( .A0(n2025), .A1(n105), .B0(n1447), .Y(n1413) );
  AOI222XLTF U734 ( .A0(n97), .A1(n174), .B0(n99), .B1(n171), .C0(n107), .C1(
        n168), .Y(n1447) );
  XOR2X1TF U735 ( .A(n1414), .B(n102), .Y(n998) );
  OAI21X1TF U736 ( .A0(n2026), .A1(n105), .B0(n1448), .Y(n1414) );
  AOI222XLTF U737 ( .A0(n97), .A1(n171), .B0(n99), .B1(n168), .C0(n107), .C1(
        n165), .Y(n1448) );
  XOR2X1TF U738 ( .A(n1415), .B(n102), .Y(n999) );
  OAI21X1TF U739 ( .A0(n2027), .A1(n105), .B0(n1449), .Y(n1415) );
  AOI222XLTF U740 ( .A0(n97), .A1(n168), .B0(n99), .B1(n165), .C0(n107), .C1(
        n162), .Y(n1449) );
  XOR2X1TF U741 ( .A(n1416), .B(n101), .Y(n1000) );
  OAI21X1TF U742 ( .A0(n2028), .A1(n105), .B0(n1450), .Y(n1416) );
  AOI222XLTF U743 ( .A0(n97), .A1(n165), .B0(n99), .B1(n162), .C0(n107), .C1(
        n159), .Y(n1450) );
  XOR2X1TF U744 ( .A(n1417), .B(n101), .Y(n1001) );
  OAI21X1TF U745 ( .A0(n2029), .A1(n105), .B0(n1451), .Y(n1417) );
  AOI222XLTF U746 ( .A0(n97), .A1(n162), .B0(n99), .B1(n159), .C0(n107), .C1(
        n156), .Y(n1451) );
  XOR2X1TF U747 ( .A(n1418), .B(n101), .Y(n1002) );
  OAI21X1TF U748 ( .A0(n2030), .A1(n104), .B0(n1452), .Y(n1418) );
  AOI222XLTF U749 ( .A0(n97), .A1(n159), .B0(n99), .B1(n156), .C0(n107), .C1(
        n153), .Y(n1452) );
  XOR2X1TF U750 ( .A(n1419), .B(n101), .Y(n1003) );
  OAI21X1TF U751 ( .A0(n2031), .A1(n104), .B0(n1453), .Y(n1419) );
  AOI222XLTF U752 ( .A0(n97), .A1(n156), .B0(n99), .B1(n153), .C0(n107), .C1(
        n150), .Y(n1453) );
  XOR2X1TF U753 ( .A(n1420), .B(n101), .Y(n1004) );
  OAI21X1TF U754 ( .A0(n2032), .A1(n104), .B0(n1454), .Y(n1420) );
  AOI222XLTF U755 ( .A0(n97), .A1(n153), .B0(n99), .B1(n150), .C0(n107), .C1(
        n147), .Y(n1454) );
  XOR2X1TF U756 ( .A(n1421), .B(n101), .Y(n1005) );
  OAI21X1TF U757 ( .A0(n2033), .A1(n104), .B0(n1455), .Y(n1421) );
  AOI222XLTF U758 ( .A0(n97), .A1(n150), .B0(n99), .B1(n147), .C0(n107), .C1(
        n144), .Y(n1455) );
  XOR2X1TF U759 ( .A(n1422), .B(n101), .Y(n1006) );
  OAI21X1TF U760 ( .A0(n2034), .A1(n104), .B0(n1456), .Y(n1422) );
  AOI222XLTF U761 ( .A0(n97), .A1(n147), .B0(n99), .B1(n144), .C0(n107), .C1(
        n141), .Y(n1456) );
  XOR2X1TF U762 ( .A(n1423), .B(n101), .Y(n1007) );
  OAI21X1TF U763 ( .A0(n2035), .A1(n104), .B0(n1457), .Y(n1423) );
  AOI222XLTF U764 ( .A0(n97), .A1(n144), .B0(n99), .B1(n141), .C0(n107), .C1(
        n138), .Y(n1457) );
  XOR2X1TF U765 ( .A(n1424), .B(n101), .Y(n1008) );
  OAI21X1TF U766 ( .A0(n2036), .A1(n104), .B0(n1458), .Y(n1424) );
  AOI222XLTF U767 ( .A0(n97), .A1(n141), .B0(n99), .B1(n138), .C0(n107), .C1(
        n135), .Y(n1458) );
  XOR2X1TF U768 ( .A(n1425), .B(n101), .Y(n1009) );
  OAI21X1TF U769 ( .A0(n2037), .A1(n104), .B0(n1459), .Y(n1425) );
  AOI222XLTF U770 ( .A0(n97), .A1(n138), .B0(n99), .B1(n135), .C0(n107), .C1(
        n132), .Y(n1459) );
  XOR2X1TF U771 ( .A(n1426), .B(n101), .Y(n1010) );
  OAI21X1TF U772 ( .A0(n104), .A1(n2038), .B0(n2298), .Y(n1426) );
  XOR2X1TF U775 ( .A(n1427), .B(n101), .Y(n1011) );
  OAI21X1TF U776 ( .A0(n104), .A1(n2039), .B0(n2309), .Y(n1427) );
  INVX2TF U779 ( .A(n91), .Y(n1012) );
  XOR2X1TF U780 ( .A(n1462), .B(n91), .Y(n1013) );
  OAI21X1TF U781 ( .A0(n2006), .A1(n94), .B0(n1496), .Y(n1462) );
  NAND2X1TF U782 ( .A(n96), .B(n225), .Y(n1496) );
  XOR2X1TF U783 ( .A(n1463), .B(n91), .Y(n1014) );
  OAI21X1TF U784 ( .A0(n2007), .A1(n94), .B0(n1497), .Y(n1463) );
  AOI21X1TF U785 ( .A0(n96), .A1(n222), .B0(n823), .Y(n1497) );
  AND2X2TF U786 ( .A(n88), .B(n225), .Y(n823) );
  XOR2X1TF U787 ( .A(n1464), .B(n91), .Y(n1015) );
  OAI21X1TF U788 ( .A0(n2008), .A1(n94), .B0(n1498), .Y(n1464) );
  AOI222XLTF U789 ( .A0(n86), .A1(n224), .B0(n88), .B1(n222), .C0(n96), .C1(
        n219), .Y(n1498) );
  XOR2X1TF U790 ( .A(n1465), .B(n91), .Y(n1016) );
  OAI21X1TF U791 ( .A0(n2009), .A1(n94), .B0(n1499), .Y(n1465) );
  AOI222XLTF U792 ( .A0(n86), .A1(n221), .B0(n88), .B1(n219), .C0(n96), .C1(
        n216), .Y(n1499) );
  XOR2X1TF U793 ( .A(n1466), .B(n91), .Y(n1017) );
  OAI21X1TF U794 ( .A0(n2010), .A1(n94), .B0(n1500), .Y(n1466) );
  AOI222XLTF U795 ( .A0(n86), .A1(n218), .B0(n88), .B1(n216), .C0(n96), .C1(
        n213), .Y(n1500) );
  XOR2X1TF U796 ( .A(n1467), .B(n91), .Y(n1018) );
  OAI21X1TF U797 ( .A0(n2011), .A1(n94), .B0(n1501), .Y(n1467) );
  AOI222XLTF U798 ( .A0(n86), .A1(n215), .B0(n88), .B1(n213), .C0(n96), .C1(
        n210), .Y(n1501) );
  XOR2X1TF U799 ( .A(n1468), .B(n91), .Y(n1019) );
  OAI21X1TF U800 ( .A0(n2012), .A1(n94), .B0(n1502), .Y(n1468) );
  AOI222XLTF U801 ( .A0(n86), .A1(n212), .B0(n88), .B1(n210), .C0(n96), .C1(
        n207), .Y(n1502) );
  XOR2X1TF U802 ( .A(n1469), .B(n91), .Y(n1020) );
  OAI21X1TF U803 ( .A0(n2013), .A1(n94), .B0(n1503), .Y(n1469) );
  AOI222XLTF U804 ( .A0(n86), .A1(n209), .B0(n88), .B1(n207), .C0(n96), .C1(
        n204), .Y(n1503) );
  XOR2X1TF U805 ( .A(n1470), .B(n91), .Y(n1021) );
  OAI21X1TF U806 ( .A0(n2014), .A1(n94), .B0(n1504), .Y(n1470) );
  AOI222XLTF U807 ( .A0(n86), .A1(n206), .B0(n88), .B1(n204), .C0(n96), .C1(
        n201), .Y(n1504) );
  XOR2X1TF U808 ( .A(n1471), .B(n91), .Y(n1022) );
  OAI21X1TF U809 ( .A0(n2015), .A1(n94), .B0(n1505), .Y(n1471) );
  AOI222XLTF U810 ( .A0(n86), .A1(n203), .B0(n88), .B1(n201), .C0(n96), .C1(
        n198), .Y(n1505) );
  XOR2X1TF U811 ( .A(n1472), .B(n90), .Y(n1023) );
  OAI21X1TF U812 ( .A0(n2016), .A1(n94), .B0(n1506), .Y(n1472) );
  AOI222XLTF U813 ( .A0(n86), .A1(n200), .B0(n88), .B1(n198), .C0(n96), .C1(
        n195), .Y(n1506) );
  XOR2X1TF U814 ( .A(n1473), .B(n90), .Y(n1024) );
  OAI21X1TF U815 ( .A0(n2017), .A1(n94), .B0(n1507), .Y(n1473) );
  AOI222XLTF U816 ( .A0(n86), .A1(n197), .B0(n88), .B1(n195), .C0(n96), .C1(
        n192), .Y(n1507) );
  XOR2X1TF U817 ( .A(n1474), .B(n90), .Y(n1025) );
  OAI21X1TF U818 ( .A0(n2018), .A1(n93), .B0(n1508), .Y(n1474) );
  AOI222XLTF U819 ( .A0(n86), .A1(n194), .B0(n88), .B1(n192), .C0(n96), .C1(
        n189), .Y(n1508) );
  XOR2X1TF U820 ( .A(n1475), .B(n90), .Y(n1026) );
  OAI21X1TF U821 ( .A0(n2019), .A1(n93), .B0(n1509), .Y(n1475) );
  AOI222XLTF U822 ( .A0(n86), .A1(n191), .B0(n88), .B1(n189), .C0(n96), .C1(
        n186), .Y(n1509) );
  XOR2X1TF U823 ( .A(n1476), .B(n90), .Y(n1027) );
  OAI21X1TF U824 ( .A0(n2020), .A1(n93), .B0(n1510), .Y(n1476) );
  AOI222XLTF U825 ( .A0(n86), .A1(n188), .B0(n88), .B1(n186), .C0(n96), .C1(
        n183), .Y(n1510) );
  XOR2X1TF U826 ( .A(n1477), .B(n90), .Y(n1028) );
  OAI21X1TF U827 ( .A0(n2021), .A1(n93), .B0(n1511), .Y(n1477) );
  AOI222XLTF U828 ( .A0(n86), .A1(n185), .B0(n88), .B1(n183), .C0(n96), .C1(
        n180), .Y(n1511) );
  XOR2X1TF U829 ( .A(n1478), .B(n90), .Y(n1029) );
  OAI21X1TF U830 ( .A0(n2022), .A1(n93), .B0(n1512), .Y(n1478) );
  AOI222XLTF U831 ( .A0(n86), .A1(n182), .B0(n88), .B1(n180), .C0(n95), .C1(
        n177), .Y(n1512) );
  XOR2X1TF U832 ( .A(n1479), .B(n90), .Y(n1030) );
  OAI21X1TF U833 ( .A0(n2023), .A1(n93), .B0(n1513), .Y(n1479) );
  AOI222XLTF U834 ( .A0(n86), .A1(n179), .B0(n87), .B1(n177), .C0(n95), .C1(
        n174), .Y(n1513) );
  XOR2X1TF U835 ( .A(n1480), .B(n90), .Y(n1031) );
  OAI21X1TF U836 ( .A0(n2024), .A1(n93), .B0(n1514), .Y(n1480) );
  AOI222XLTF U837 ( .A0(n85), .A1(n176), .B0(n87), .B1(n174), .C0(n95), .C1(
        n171), .Y(n1514) );
  XOR2X1TF U838 ( .A(n1481), .B(n90), .Y(n1032) );
  OAI21X1TF U839 ( .A0(n2025), .A1(n93), .B0(n1515), .Y(n1481) );
  AOI222XLTF U840 ( .A0(n85), .A1(n173), .B0(n87), .B1(n171), .C0(n95), .C1(
        n168), .Y(n1515) );
  XOR2X1TF U841 ( .A(n1482), .B(n90), .Y(n1033) );
  OAI21X1TF U842 ( .A0(n2026), .A1(n93), .B0(n1516), .Y(n1482) );
  AOI222XLTF U843 ( .A0(n85), .A1(n170), .B0(n87), .B1(n168), .C0(n95), .C1(
        n165), .Y(n1516) );
  XOR2X1TF U844 ( .A(n1483), .B(n90), .Y(n1034) );
  OAI21X1TF U845 ( .A0(n2027), .A1(n93), .B0(n1517), .Y(n1483) );
  AOI222XLTF U846 ( .A0(n85), .A1(n167), .B0(n87), .B1(n165), .C0(n95), .C1(
        n162), .Y(n1517) );
  XOR2X1TF U847 ( .A(n1484), .B(n89), .Y(n1035) );
  OAI21X1TF U848 ( .A0(n2028), .A1(n93), .B0(n1518), .Y(n1484) );
  AOI222XLTF U849 ( .A0(n85), .A1(n164), .B0(n87), .B1(n162), .C0(n95), .C1(
        n159), .Y(n1518) );
  XOR2X1TF U850 ( .A(n1485), .B(n89), .Y(n1036) );
  OAI21X1TF U851 ( .A0(n2029), .A1(n93), .B0(n1519), .Y(n1485) );
  AOI222XLTF U852 ( .A0(n85), .A1(n161), .B0(n87), .B1(n159), .C0(n95), .C1(
        n156), .Y(n1519) );
  XOR2X1TF U853 ( .A(n1486), .B(n89), .Y(n1037) );
  OAI21X1TF U854 ( .A0(n2030), .A1(n92), .B0(n1520), .Y(n1486) );
  AOI222XLTF U855 ( .A0(n85), .A1(n158), .B0(n87), .B1(n156), .C0(n95), .C1(
        n153), .Y(n1520) );
  XOR2X1TF U856 ( .A(n1487), .B(n89), .Y(n1038) );
  OAI21X1TF U857 ( .A0(n2031), .A1(n92), .B0(n1521), .Y(n1487) );
  AOI222XLTF U858 ( .A0(n85), .A1(n155), .B0(n87), .B1(n153), .C0(n95), .C1(
        n150), .Y(n1521) );
  XOR2X1TF U859 ( .A(n1488), .B(n89), .Y(n1039) );
  OAI21X1TF U860 ( .A0(n2032), .A1(n92), .B0(n1522), .Y(n1488) );
  AOI222XLTF U861 ( .A0(n85), .A1(n152), .B0(n87), .B1(n150), .C0(n95), .C1(
        n147), .Y(n1522) );
  XOR2X1TF U862 ( .A(n1489), .B(n89), .Y(n1040) );
  OAI21X1TF U863 ( .A0(n2033), .A1(n92), .B0(n1523), .Y(n1489) );
  AOI222XLTF U864 ( .A0(n85), .A1(n149), .B0(n87), .B1(n147), .C0(n95), .C1(
        n144), .Y(n1523) );
  XOR2X1TF U865 ( .A(n1490), .B(n89), .Y(n1041) );
  OAI21X1TF U866 ( .A0(n2034), .A1(n92), .B0(n1524), .Y(n1490) );
  AOI222XLTF U867 ( .A0(n85), .A1(n146), .B0(n87), .B1(n144), .C0(n95), .C1(
        n141), .Y(n1524) );
  XOR2X1TF U868 ( .A(n1491), .B(n89), .Y(n1042) );
  OAI21X1TF U869 ( .A0(n2035), .A1(n92), .B0(n1525), .Y(n1491) );
  AOI222XLTF U870 ( .A0(n85), .A1(n143), .B0(n87), .B1(n141), .C0(n95), .C1(
        n138), .Y(n1525) );
  XOR2X1TF U871 ( .A(n1492), .B(n89), .Y(n1043) );
  OAI21X1TF U872 ( .A0(n2036), .A1(n92), .B0(n1526), .Y(n1492) );
  AOI222XLTF U873 ( .A0(n85), .A1(n140), .B0(n87), .B1(n138), .C0(n95), .C1(
        n135), .Y(n1526) );
  XOR2X1TF U874 ( .A(n1493), .B(n89), .Y(n1044) );
  OAI21X1TF U875 ( .A0(n2037), .A1(n92), .B0(n1527), .Y(n1493) );
  AOI222XLTF U876 ( .A0(n85), .A1(n137), .B0(n87), .B1(n135), .C0(n95), .C1(
        n132), .Y(n1527) );
  XOR2X1TF U877 ( .A(n1494), .B(n89), .Y(n1045) );
  OAI21X1TF U878 ( .A0(n92), .A1(n2038), .B0(n2297), .Y(n1494) );
  XOR2X1TF U881 ( .A(n1495), .B(n89), .Y(n1046) );
  OAI21X1TF U882 ( .A0(n92), .A1(n2039), .B0(n2308), .Y(n1495) );
  INVX2TF U885 ( .A(n79), .Y(n1047) );
  XOR2X1TF U886 ( .A(n1530), .B(n79), .Y(n1048) );
  OAI21X1TF U887 ( .A0(n2006), .A1(n82), .B0(n1564), .Y(n1530) );
  NAND2X1TF U888 ( .A(n84), .B(n224), .Y(n1564) );
  XOR2X1TF U889 ( .A(n1531), .B(n79), .Y(n1049) );
  OAI21X1TF U890 ( .A0(n2007), .A1(n82), .B0(n1565), .Y(n1531) );
  AOI21X1TF U891 ( .A0(n84), .A1(n221), .B0(n826), .Y(n1565) );
  AND2X2TF U892 ( .A(n76), .B(n224), .Y(n826) );
  XOR2X1TF U893 ( .A(n1532), .B(n79), .Y(n1050) );
  OAI21X1TF U894 ( .A0(n2008), .A1(n82), .B0(n1566), .Y(n1532) );
  AOI222XLTF U895 ( .A0(n74), .A1(n224), .B0(n76), .B1(n221), .C0(n84), .C1(
        n218), .Y(n1566) );
  XOR2X1TF U896 ( .A(n1533), .B(n79), .Y(n1051) );
  OAI21X1TF U897 ( .A0(n2009), .A1(n82), .B0(n1567), .Y(n1533) );
  AOI222XLTF U898 ( .A0(n74), .A1(n221), .B0(n76), .B1(n218), .C0(n84), .C1(
        n215), .Y(n1567) );
  XOR2X1TF U899 ( .A(n1534), .B(n79), .Y(n1052) );
  OAI21X1TF U900 ( .A0(n2010), .A1(n82), .B0(n1568), .Y(n1534) );
  AOI222XLTF U901 ( .A0(n74), .A1(n218), .B0(n76), .B1(n215), .C0(n84), .C1(
        n212), .Y(n1568) );
  XOR2X1TF U902 ( .A(n1535), .B(n79), .Y(n1053) );
  OAI21X1TF U903 ( .A0(n2011), .A1(n82), .B0(n1569), .Y(n1535) );
  AOI222XLTF U904 ( .A0(n74), .A1(n215), .B0(n76), .B1(n212), .C0(n84), .C1(
        n209), .Y(n1569) );
  XOR2X1TF U905 ( .A(n1536), .B(n79), .Y(n1054) );
  OAI21X1TF U906 ( .A0(n2012), .A1(n82), .B0(n1570), .Y(n1536) );
  AOI222XLTF U907 ( .A0(n74), .A1(n212), .B0(n76), .B1(n209), .C0(n84), .C1(
        n206), .Y(n1570) );
  XOR2X1TF U908 ( .A(n1537), .B(n79), .Y(n1055) );
  OAI21X1TF U909 ( .A0(n2013), .A1(n82), .B0(n1571), .Y(n1537) );
  AOI222XLTF U910 ( .A0(n74), .A1(n209), .B0(n76), .B1(n206), .C0(n84), .C1(
        n203), .Y(n1571) );
  XOR2X1TF U911 ( .A(n1538), .B(n79), .Y(n1056) );
  OAI21X1TF U912 ( .A0(n2014), .A1(n82), .B0(n1572), .Y(n1538) );
  AOI222XLTF U913 ( .A0(n74), .A1(n206), .B0(n76), .B1(n203), .C0(n84), .C1(
        n200), .Y(n1572) );
  XOR2X1TF U914 ( .A(n1539), .B(n79), .Y(n1057) );
  OAI21X1TF U915 ( .A0(n2015), .A1(n82), .B0(n1573), .Y(n1539) );
  AOI222XLTF U916 ( .A0(n74), .A1(n203), .B0(n76), .B1(n200), .C0(n84), .C1(
        n197), .Y(n1573) );
  XOR2X1TF U917 ( .A(n1540), .B(n78), .Y(n1058) );
  OAI21X1TF U918 ( .A0(n2016), .A1(n82), .B0(n1574), .Y(n1540) );
  AOI222XLTF U919 ( .A0(n74), .A1(n200), .B0(n76), .B1(n197), .C0(n84), .C1(
        n194), .Y(n1574) );
  XOR2X1TF U920 ( .A(n1541), .B(n78), .Y(n1059) );
  OAI21X1TF U921 ( .A0(n2017), .A1(n82), .B0(n1575), .Y(n1541) );
  AOI222XLTF U922 ( .A0(n74), .A1(n197), .B0(n76), .B1(n194), .C0(n84), .C1(
        n191), .Y(n1575) );
  XOR2X1TF U923 ( .A(n1542), .B(n78), .Y(n1060) );
  OAI21X1TF U924 ( .A0(n2018), .A1(n81), .B0(n1576), .Y(n1542) );
  AOI222XLTF U925 ( .A0(n74), .A1(n194), .B0(n76), .B1(n191), .C0(n84), .C1(
        n188), .Y(n1576) );
  XOR2X1TF U926 ( .A(n1543), .B(n78), .Y(n1061) );
  OAI21X1TF U927 ( .A0(n2019), .A1(n81), .B0(n1577), .Y(n1543) );
  AOI222XLTF U928 ( .A0(n74), .A1(n191), .B0(n76), .B1(n188), .C0(n84), .C1(
        n185), .Y(n1577) );
  XOR2X1TF U929 ( .A(n1544), .B(n78), .Y(n1062) );
  OAI21X1TF U930 ( .A0(n2020), .A1(n81), .B0(n1578), .Y(n1544) );
  AOI222XLTF U931 ( .A0(n74), .A1(n188), .B0(n76), .B1(n185), .C0(n84), .C1(
        n182), .Y(n1578) );
  XOR2X1TF U932 ( .A(n1545), .B(n78), .Y(n1063) );
  OAI21X1TF U933 ( .A0(n2021), .A1(n81), .B0(n1579), .Y(n1545) );
  AOI222XLTF U934 ( .A0(n74), .A1(n185), .B0(n76), .B1(n182), .C0(n84), .C1(
        n179), .Y(n1579) );
  XOR2X1TF U935 ( .A(n1546), .B(n78), .Y(n1064) );
  OAI21X1TF U936 ( .A0(n2022), .A1(n81), .B0(n1580), .Y(n1546) );
  AOI222XLTF U937 ( .A0(n74), .A1(n182), .B0(n76), .B1(n179), .C0(n83), .C1(
        n176), .Y(n1580) );
  XOR2X1TF U938 ( .A(n1547), .B(n78), .Y(n1065) );
  OAI21X1TF U939 ( .A0(n2023), .A1(n81), .B0(n1581), .Y(n1547) );
  AOI222XLTF U940 ( .A0(n74), .A1(n179), .B0(n75), .B1(n176), .C0(n83), .C1(
        n173), .Y(n1581) );
  XOR2X1TF U941 ( .A(n1548), .B(n78), .Y(n1066) );
  OAI21X1TF U942 ( .A0(n2024), .A1(n81), .B0(n1582), .Y(n1548) );
  AOI222XLTF U943 ( .A0(n73), .A1(n176), .B0(n75), .B1(n173), .C0(n83), .C1(
        n170), .Y(n1582) );
  XOR2X1TF U944 ( .A(n1549), .B(n78), .Y(n1067) );
  OAI21X1TF U945 ( .A0(n2025), .A1(n81), .B0(n1583), .Y(n1549) );
  AOI222XLTF U946 ( .A0(n73), .A1(n173), .B0(n75), .B1(n170), .C0(n83), .C1(
        n167), .Y(n1583) );
  XOR2X1TF U947 ( .A(n1550), .B(n78), .Y(n1068) );
  OAI21X1TF U948 ( .A0(n2026), .A1(n81), .B0(n1584), .Y(n1550) );
  AOI222XLTF U949 ( .A0(n73), .A1(n170), .B0(n75), .B1(n167), .C0(n83), .C1(
        n164), .Y(n1584) );
  XOR2X1TF U950 ( .A(n1551), .B(n78), .Y(n1069) );
  OAI21X1TF U951 ( .A0(n2027), .A1(n81), .B0(n1585), .Y(n1551) );
  AOI222XLTF U952 ( .A0(n73), .A1(n167), .B0(n75), .B1(n164), .C0(n83), .C1(
        n161), .Y(n1585) );
  XOR2X1TF U953 ( .A(n1552), .B(n77), .Y(n1070) );
  OAI21X1TF U954 ( .A0(n2028), .A1(n81), .B0(n1586), .Y(n1552) );
  AOI222XLTF U955 ( .A0(n73), .A1(n164), .B0(n75), .B1(n161), .C0(n83), .C1(
        n158), .Y(n1586) );
  XOR2X1TF U956 ( .A(n1553), .B(n77), .Y(n1071) );
  OAI21X1TF U957 ( .A0(n2029), .A1(n81), .B0(n1587), .Y(n1553) );
  AOI222XLTF U958 ( .A0(n73), .A1(n161), .B0(n75), .B1(n158), .C0(n83), .C1(
        n155), .Y(n1587) );
  XOR2X1TF U959 ( .A(n1554), .B(n77), .Y(n1072) );
  OAI21X1TF U960 ( .A0(n2030), .A1(n80), .B0(n1588), .Y(n1554) );
  AOI222XLTF U961 ( .A0(n73), .A1(n158), .B0(n75), .B1(n155), .C0(n83), .C1(
        n152), .Y(n1588) );
  XOR2X1TF U962 ( .A(n1555), .B(n77), .Y(n1073) );
  OAI21X1TF U963 ( .A0(n2031), .A1(n80), .B0(n1589), .Y(n1555) );
  AOI222XLTF U964 ( .A0(n73), .A1(n155), .B0(n75), .B1(n152), .C0(n83), .C1(
        n149), .Y(n1589) );
  XOR2X1TF U965 ( .A(n1556), .B(n77), .Y(n1074) );
  OAI21X1TF U966 ( .A0(n2032), .A1(n80), .B0(n1590), .Y(n1556) );
  AOI222XLTF U967 ( .A0(n73), .A1(n152), .B0(n75), .B1(n149), .C0(n83), .C1(
        n146), .Y(n1590) );
  XOR2X1TF U968 ( .A(n1557), .B(n77), .Y(n1075) );
  OAI21X1TF U969 ( .A0(n2033), .A1(n80), .B0(n1591), .Y(n1557) );
  AOI222XLTF U970 ( .A0(n73), .A1(n149), .B0(n75), .B1(n146), .C0(n83), .C1(
        n143), .Y(n1591) );
  XOR2X1TF U971 ( .A(n1558), .B(n77), .Y(n1076) );
  OAI21X1TF U972 ( .A0(n2034), .A1(n80), .B0(n1592), .Y(n1558) );
  AOI222XLTF U973 ( .A0(n73), .A1(n146), .B0(n75), .B1(n143), .C0(n83), .C1(
        n140), .Y(n1592) );
  XOR2X1TF U974 ( .A(n1559), .B(n77), .Y(n1077) );
  OAI21X1TF U975 ( .A0(n2035), .A1(n80), .B0(n1593), .Y(n1559) );
  AOI222XLTF U976 ( .A0(n73), .A1(n143), .B0(n75), .B1(n140), .C0(n83), .C1(
        n137), .Y(n1593) );
  XOR2X1TF U977 ( .A(n1560), .B(n77), .Y(n1078) );
  OAI21X1TF U978 ( .A0(n2036), .A1(n80), .B0(n1594), .Y(n1560) );
  AOI222XLTF U979 ( .A0(n73), .A1(n140), .B0(n75), .B1(n137), .C0(n83), .C1(
        n134), .Y(n1594) );
  XOR2X1TF U980 ( .A(n1561), .B(n77), .Y(n1079) );
  OAI21X1TF U981 ( .A0(n2037), .A1(n80), .B0(n1595), .Y(n1561) );
  AOI222XLTF U982 ( .A0(n73), .A1(n137), .B0(n75), .B1(n134), .C0(n83), .C1(
        n131), .Y(n1595) );
  XOR2X1TF U983 ( .A(n1562), .B(n77), .Y(n1080) );
  OAI21X1TF U984 ( .A0(n80), .A1(n2038), .B0(n2296), .Y(n1562) );
  XOR2X1TF U987 ( .A(n1563), .B(n77), .Y(n1081) );
  OAI21X1TF U988 ( .A0(n80), .A1(n2039), .B0(n2307), .Y(n1563) );
  INVX2TF U991 ( .A(n67), .Y(n1082) );
  XOR2X1TF U992 ( .A(n1598), .B(n67), .Y(n1083) );
  OAI21X1TF U993 ( .A0(n2006), .A1(n70), .B0(n1632), .Y(n1598) );
  NAND2X1TF U994 ( .A(n72), .B(n224), .Y(n1632) );
  XOR2X1TF U995 ( .A(n1599), .B(n67), .Y(n1084) );
  OAI21X1TF U996 ( .A0(n2007), .A1(n70), .B0(n1633), .Y(n1599) );
  AOI21X1TF U997 ( .A0(n72), .A1(n221), .B0(n829), .Y(n1633) );
  AND2X2TF U998 ( .A(n64), .B(n224), .Y(n829) );
  XOR2X1TF U999 ( .A(n1600), .B(n67), .Y(n1085) );
  OAI21X1TF U1000 ( .A0(n2008), .A1(n70), .B0(n1634), .Y(n1600) );
  AOI222XLTF U1001 ( .A0(n62), .A1(n224), .B0(n64), .B1(n221), .C0(n72), .C1(
        n218), .Y(n1634) );
  XOR2X1TF U1002 ( .A(n1601), .B(n67), .Y(n1086) );
  OAI21X1TF U1003 ( .A0(n2009), .A1(n70), .B0(n1635), .Y(n1601) );
  AOI222XLTF U1004 ( .A0(n62), .A1(n221), .B0(n64), .B1(n218), .C0(n72), .C1(
        n215), .Y(n1635) );
  XOR2X1TF U1005 ( .A(n1602), .B(n67), .Y(n1087) );
  OAI21X1TF U1006 ( .A0(n2010), .A1(n70), .B0(n1636), .Y(n1602) );
  AOI222XLTF U1007 ( .A0(n62), .A1(n218), .B0(n64), .B1(n215), .C0(n72), .C1(
        n212), .Y(n1636) );
  XOR2X1TF U1008 ( .A(n1603), .B(n67), .Y(n1088) );
  OAI21X1TF U1009 ( .A0(n2011), .A1(n70), .B0(n1637), .Y(n1603) );
  AOI222XLTF U1010 ( .A0(n62), .A1(n215), .B0(n64), .B1(n212), .C0(n72), .C1(
        n209), .Y(n1637) );
  XOR2X1TF U1011 ( .A(n1604), .B(n67), .Y(n1089) );
  OAI21X1TF U1012 ( .A0(n2012), .A1(n70), .B0(n1638), .Y(n1604) );
  AOI222XLTF U1013 ( .A0(n62), .A1(n212), .B0(n64), .B1(n209), .C0(n72), .C1(
        n206), .Y(n1638) );
  XOR2X1TF U1014 ( .A(n1605), .B(n67), .Y(n1090) );
  OAI21X1TF U1015 ( .A0(n2013), .A1(n70), .B0(n1639), .Y(n1605) );
  AOI222XLTF U1016 ( .A0(n62), .A1(n209), .B0(n64), .B1(n206), .C0(n72), .C1(
        n203), .Y(n1639) );
  XOR2X1TF U1017 ( .A(n1606), .B(n67), .Y(n1091) );
  OAI21X1TF U1018 ( .A0(n2014), .A1(n70), .B0(n1640), .Y(n1606) );
  AOI222XLTF U1019 ( .A0(n62), .A1(n206), .B0(n64), .B1(n203), .C0(n72), .C1(
        n200), .Y(n1640) );
  XOR2X1TF U1020 ( .A(n1607), .B(n67), .Y(n1092) );
  OAI21X1TF U1021 ( .A0(n2015), .A1(n70), .B0(n1641), .Y(n1607) );
  AOI222XLTF U1022 ( .A0(n62), .A1(n203), .B0(n64), .B1(n200), .C0(n72), .C1(
        n197), .Y(n1641) );
  XOR2X1TF U1023 ( .A(n1608), .B(n66), .Y(n1093) );
  OAI21X1TF U1024 ( .A0(n2016), .A1(n70), .B0(n1642), .Y(n1608) );
  AOI222XLTF U1025 ( .A0(n62), .A1(n200), .B0(n64), .B1(n197), .C0(n72), .C1(
        n194), .Y(n1642) );
  XOR2X1TF U1026 ( .A(n1609), .B(n66), .Y(n1094) );
  OAI21X1TF U1027 ( .A0(n2017), .A1(n70), .B0(n1643), .Y(n1609) );
  AOI222XLTF U1028 ( .A0(n62), .A1(n197), .B0(n64), .B1(n194), .C0(n72), .C1(
        n191), .Y(n1643) );
  XOR2X1TF U1029 ( .A(n1610), .B(n66), .Y(n1095) );
  OAI21X1TF U1030 ( .A0(n2018), .A1(n69), .B0(n1644), .Y(n1610) );
  AOI222XLTF U1031 ( .A0(n62), .A1(n194), .B0(n64), .B1(n191), .C0(n72), .C1(
        n188), .Y(n1644) );
  XOR2X1TF U1032 ( .A(n1611), .B(n66), .Y(n1096) );
  OAI21X1TF U1033 ( .A0(n2019), .A1(n69), .B0(n1645), .Y(n1611) );
  AOI222XLTF U1034 ( .A0(n62), .A1(n191), .B0(n64), .B1(n188), .C0(n72), .C1(
        n185), .Y(n1645) );
  XOR2X1TF U1035 ( .A(n1612), .B(n66), .Y(n1097) );
  OAI21X1TF U1036 ( .A0(n2020), .A1(n69), .B0(n1646), .Y(n1612) );
  AOI222XLTF U1037 ( .A0(n62), .A1(n188), .B0(n64), .B1(n185), .C0(n72), .C1(
        n182), .Y(n1646) );
  XOR2X1TF U1038 ( .A(n1613), .B(n66), .Y(n1098) );
  OAI21X1TF U1039 ( .A0(n2021), .A1(n69), .B0(n1647), .Y(n1613) );
  AOI222XLTF U1040 ( .A0(n62), .A1(n185), .B0(n64), .B1(n182), .C0(n72), .C1(
        n179), .Y(n1647) );
  XOR2X1TF U1041 ( .A(n1614), .B(n66), .Y(n1099) );
  OAI21X1TF U1042 ( .A0(n2022), .A1(n69), .B0(n1648), .Y(n1614) );
  AOI222XLTF U1043 ( .A0(n62), .A1(n182), .B0(n64), .B1(n179), .C0(n71), .C1(
        n176), .Y(n1648) );
  XOR2X1TF U1044 ( .A(n1615), .B(n66), .Y(n1100) );
  OAI21X1TF U1045 ( .A0(n2023), .A1(n69), .B0(n1649), .Y(n1615) );
  AOI222XLTF U1046 ( .A0(n62), .A1(n179), .B0(n63), .B1(n176), .C0(n71), .C1(
        n173), .Y(n1649) );
  XOR2X1TF U1047 ( .A(n1616), .B(n66), .Y(n1101) );
  OAI21X1TF U1048 ( .A0(n2024), .A1(n69), .B0(n1650), .Y(n1616) );
  AOI222XLTF U1049 ( .A0(n61), .A1(n176), .B0(n63), .B1(n173), .C0(n71), .C1(
        n170), .Y(n1650) );
  XOR2X1TF U1050 ( .A(n1617), .B(n66), .Y(n1102) );
  OAI21X1TF U1051 ( .A0(n2025), .A1(n69), .B0(n1651), .Y(n1617) );
  AOI222XLTF U1052 ( .A0(n61), .A1(n173), .B0(n63), .B1(n170), .C0(n71), .C1(
        n167), .Y(n1651) );
  XOR2X1TF U1053 ( .A(n1618), .B(n66), .Y(n1103) );
  OAI21X1TF U1054 ( .A0(n2026), .A1(n69), .B0(n1652), .Y(n1618) );
  AOI222XLTF U1055 ( .A0(n61), .A1(n170), .B0(n63), .B1(n167), .C0(n71), .C1(
        n164), .Y(n1652) );
  XOR2X1TF U1056 ( .A(n1619), .B(n66), .Y(n1104) );
  OAI21X1TF U1057 ( .A0(n2027), .A1(n69), .B0(n1653), .Y(n1619) );
  AOI222XLTF U1058 ( .A0(n61), .A1(n167), .B0(n63), .B1(n164), .C0(n71), .C1(
        n161), .Y(n1653) );
  XOR2X1TF U1059 ( .A(n1620), .B(n65), .Y(n1105) );
  OAI21X1TF U1060 ( .A0(n2028), .A1(n69), .B0(n1654), .Y(n1620) );
  AOI222XLTF U1061 ( .A0(n61), .A1(n164), .B0(n63), .B1(n161), .C0(n71), .C1(
        n158), .Y(n1654) );
  XOR2X1TF U1062 ( .A(n1621), .B(n65), .Y(n1106) );
  OAI21X1TF U1063 ( .A0(n2029), .A1(n69), .B0(n1655), .Y(n1621) );
  AOI222XLTF U1064 ( .A0(n61), .A1(n161), .B0(n63), .B1(n158), .C0(n71), .C1(
        n155), .Y(n1655) );
  XOR2X1TF U1065 ( .A(n1622), .B(n65), .Y(n1107) );
  OAI21X1TF U1066 ( .A0(n2030), .A1(n68), .B0(n1656), .Y(n1622) );
  AOI222XLTF U1067 ( .A0(n61), .A1(n158), .B0(n63), .B1(n155), .C0(n71), .C1(
        n152), .Y(n1656) );
  XOR2X1TF U1068 ( .A(n1623), .B(n65), .Y(n1108) );
  OAI21X1TF U1069 ( .A0(n2031), .A1(n68), .B0(n1657), .Y(n1623) );
  AOI222XLTF U1070 ( .A0(n61), .A1(n155), .B0(n63), .B1(n152), .C0(n71), .C1(
        n149), .Y(n1657) );
  XOR2X1TF U1071 ( .A(n1624), .B(n65), .Y(n1109) );
  OAI21X1TF U1072 ( .A0(n2032), .A1(n68), .B0(n1658), .Y(n1624) );
  AOI222XLTF U1073 ( .A0(n61), .A1(n152), .B0(n63), .B1(n149), .C0(n71), .C1(
        n146), .Y(n1658) );
  XOR2X1TF U1074 ( .A(n1625), .B(n65), .Y(n1110) );
  OAI21X1TF U1075 ( .A0(n2033), .A1(n68), .B0(n1659), .Y(n1625) );
  AOI222XLTF U1076 ( .A0(n61), .A1(n149), .B0(n63), .B1(n146), .C0(n71), .C1(
        n143), .Y(n1659) );
  XOR2X1TF U1077 ( .A(n1626), .B(n65), .Y(n1111) );
  OAI21X1TF U1078 ( .A0(n2034), .A1(n68), .B0(n1660), .Y(n1626) );
  AOI222XLTF U1079 ( .A0(n61), .A1(n146), .B0(n63), .B1(n143), .C0(n71), .C1(
        n140), .Y(n1660) );
  XOR2X1TF U1080 ( .A(n1627), .B(n65), .Y(n1112) );
  OAI21X1TF U1081 ( .A0(n2035), .A1(n68), .B0(n1661), .Y(n1627) );
  AOI222XLTF U1082 ( .A0(n61), .A1(n143), .B0(n63), .B1(n140), .C0(n71), .C1(
        n137), .Y(n1661) );
  XOR2X1TF U1083 ( .A(n1628), .B(n65), .Y(n1113) );
  OAI21X1TF U1084 ( .A0(n2036), .A1(n68), .B0(n1662), .Y(n1628) );
  AOI222XLTF U1085 ( .A0(n61), .A1(n140), .B0(n63), .B1(n137), .C0(n71), .C1(
        n134), .Y(n1662) );
  XOR2X1TF U1086 ( .A(n1629), .B(n65), .Y(n1114) );
  OAI21X1TF U1087 ( .A0(n2037), .A1(n68), .B0(n1663), .Y(n1629) );
  AOI222XLTF U1088 ( .A0(n61), .A1(n137), .B0(n63), .B1(n134), .C0(n71), .C1(
        n131), .Y(n1663) );
  XOR2X1TF U1089 ( .A(n1630), .B(n65), .Y(n1115) );
  OAI21X1TF U1090 ( .A0(n68), .A1(n2038), .B0(n2295), .Y(n1630) );
  XOR2X1TF U1093 ( .A(n1631), .B(n65), .Y(n1116) );
  OAI21X1TF U1094 ( .A0(n68), .A1(n2039), .B0(n2306), .Y(n1631) );
  INVX2TF U1097 ( .A(n55), .Y(n1117) );
  XOR2X1TF U1098 ( .A(n1666), .B(n55), .Y(n1118) );
  OAI21X1TF U1099 ( .A0(n2006), .A1(n58), .B0(n1700), .Y(n1666) );
  NAND2X1TF U1100 ( .A(n60), .B(n224), .Y(n1700) );
  XOR2X1TF U1101 ( .A(n1667), .B(n55), .Y(n1119) );
  OAI21X1TF U1102 ( .A0(n2007), .A1(n58), .B0(n1701), .Y(n1667) );
  AOI21X1TF U1103 ( .A0(n60), .A1(n221), .B0(n832), .Y(n1701) );
  AND2X2TF U1104 ( .A(n52), .B(n224), .Y(n832) );
  XOR2X1TF U1105 ( .A(n1668), .B(n55), .Y(n1120) );
  OAI21X1TF U1106 ( .A0(n2008), .A1(n58), .B0(n1702), .Y(n1668) );
  AOI222XLTF U1107 ( .A0(n50), .A1(n224), .B0(n52), .B1(n221), .C0(n60), .C1(
        n218), .Y(n1702) );
  XOR2X1TF U1108 ( .A(n1669), .B(n55), .Y(n1121) );
  OAI21X1TF U1109 ( .A0(n2009), .A1(n58), .B0(n1703), .Y(n1669) );
  AOI222XLTF U1110 ( .A0(n50), .A1(n221), .B0(n52), .B1(n218), .C0(n60), .C1(
        n215), .Y(n1703) );
  XOR2X1TF U1111 ( .A(n1670), .B(n55), .Y(n1122) );
  OAI21X1TF U1112 ( .A0(n2010), .A1(n58), .B0(n1704), .Y(n1670) );
  AOI222XLTF U1113 ( .A0(n50), .A1(n218), .B0(n52), .B1(n215), .C0(n60), .C1(
        n212), .Y(n1704) );
  XOR2X1TF U1114 ( .A(n1671), .B(n55), .Y(n1123) );
  OAI21X1TF U1115 ( .A0(n2011), .A1(n58), .B0(n1705), .Y(n1671) );
  AOI222XLTF U1116 ( .A0(n50), .A1(n215), .B0(n52), .B1(n212), .C0(n60), .C1(
        n209), .Y(n1705) );
  XOR2X1TF U1117 ( .A(n1672), .B(n55), .Y(n1124) );
  OAI21X1TF U1118 ( .A0(n2012), .A1(n58), .B0(n1706), .Y(n1672) );
  AOI222XLTF U1119 ( .A0(n50), .A1(n212), .B0(n52), .B1(n209), .C0(n60), .C1(
        n206), .Y(n1706) );
  XOR2X1TF U1120 ( .A(n1673), .B(n55), .Y(n1125) );
  OAI21X1TF U1121 ( .A0(n2013), .A1(n58), .B0(n1707), .Y(n1673) );
  AOI222XLTF U1122 ( .A0(n50), .A1(n209), .B0(n52), .B1(n206), .C0(n60), .C1(
        n203), .Y(n1707) );
  XOR2X1TF U1123 ( .A(n1674), .B(n55), .Y(n1126) );
  OAI21X1TF U1124 ( .A0(n2014), .A1(n58), .B0(n1708), .Y(n1674) );
  AOI222XLTF U1125 ( .A0(n50), .A1(n206), .B0(n52), .B1(n203), .C0(n60), .C1(
        n200), .Y(n1708) );
  XOR2X1TF U1126 ( .A(n1675), .B(n55), .Y(n1127) );
  OAI21X1TF U1127 ( .A0(n2015), .A1(n58), .B0(n1709), .Y(n1675) );
  AOI222XLTF U1128 ( .A0(n50), .A1(n203), .B0(n52), .B1(n200), .C0(n60), .C1(
        n197), .Y(n1709) );
  XOR2X1TF U1129 ( .A(n1676), .B(n54), .Y(n1128) );
  OAI21X1TF U1130 ( .A0(n2016), .A1(n58), .B0(n1710), .Y(n1676) );
  AOI222XLTF U1131 ( .A0(n50), .A1(n200), .B0(n52), .B1(n197), .C0(n60), .C1(
        n194), .Y(n1710) );
  XOR2X1TF U1132 ( .A(n1677), .B(n54), .Y(n1129) );
  OAI21X1TF U1133 ( .A0(n2017), .A1(n58), .B0(n1711), .Y(n1677) );
  AOI222XLTF U1134 ( .A0(n50), .A1(n197), .B0(n52), .B1(n194), .C0(n60), .C1(
        n191), .Y(n1711) );
  XOR2X1TF U1135 ( .A(n1678), .B(n54), .Y(n1130) );
  OAI21X1TF U1136 ( .A0(n2018), .A1(n57), .B0(n1712), .Y(n1678) );
  AOI222XLTF U1137 ( .A0(n50), .A1(n194), .B0(n52), .B1(n191), .C0(n60), .C1(
        n188), .Y(n1712) );
  XOR2X1TF U1138 ( .A(n1679), .B(n54), .Y(n1131) );
  OAI21X1TF U1139 ( .A0(n2019), .A1(n57), .B0(n1713), .Y(n1679) );
  AOI222XLTF U1140 ( .A0(n50), .A1(n191), .B0(n52), .B1(n188), .C0(n60), .C1(
        n185), .Y(n1713) );
  XOR2X1TF U1141 ( .A(n1680), .B(n54), .Y(n1132) );
  OAI21X1TF U1142 ( .A0(n2020), .A1(n57), .B0(n1714), .Y(n1680) );
  AOI222XLTF U1143 ( .A0(n50), .A1(n188), .B0(n52), .B1(n185), .C0(n60), .C1(
        n182), .Y(n1714) );
  XOR2X1TF U1144 ( .A(n1681), .B(n54), .Y(n1133) );
  OAI21X1TF U1145 ( .A0(n2021), .A1(n57), .B0(n1715), .Y(n1681) );
  AOI222XLTF U1146 ( .A0(n50), .A1(n185), .B0(n52), .B1(n182), .C0(n60), .C1(
        n179), .Y(n1715) );
  XOR2X1TF U1147 ( .A(n1682), .B(n54), .Y(n1134) );
  OAI21X1TF U1148 ( .A0(n2022), .A1(n57), .B0(n1716), .Y(n1682) );
  AOI222XLTF U1149 ( .A0(n50), .A1(n182), .B0(n52), .B1(n179), .C0(n59), .C1(
        n176), .Y(n1716) );
  XOR2X1TF U1150 ( .A(n1683), .B(n54), .Y(n1135) );
  OAI21X1TF U1151 ( .A0(n2023), .A1(n57), .B0(n1717), .Y(n1683) );
  AOI222XLTF U1152 ( .A0(n50), .A1(n179), .B0(n51), .B1(n176), .C0(n59), .C1(
        n173), .Y(n1717) );
  XOR2X1TF U1153 ( .A(n1684), .B(n54), .Y(n1136) );
  OAI21X1TF U1154 ( .A0(n2024), .A1(n57), .B0(n1718), .Y(n1684) );
  AOI222XLTF U1155 ( .A0(n49), .A1(n176), .B0(n51), .B1(n173), .C0(n59), .C1(
        n170), .Y(n1718) );
  XOR2X1TF U1156 ( .A(n1685), .B(n54), .Y(n1137) );
  OAI21X1TF U1157 ( .A0(n2025), .A1(n57), .B0(n1719), .Y(n1685) );
  AOI222XLTF U1158 ( .A0(n49), .A1(n173), .B0(n51), .B1(n170), .C0(n59), .C1(
        n167), .Y(n1719) );
  XOR2X1TF U1159 ( .A(n1686), .B(n54), .Y(n1138) );
  OAI21X1TF U1160 ( .A0(n2026), .A1(n57), .B0(n1720), .Y(n1686) );
  AOI222XLTF U1161 ( .A0(n49), .A1(n170), .B0(n51), .B1(n167), .C0(n59), .C1(
        n164), .Y(n1720) );
  XOR2X1TF U1162 ( .A(n1687), .B(n54), .Y(n1139) );
  OAI21X1TF U1163 ( .A0(n2027), .A1(n57), .B0(n1721), .Y(n1687) );
  AOI222XLTF U1164 ( .A0(n49), .A1(n167), .B0(n51), .B1(n164), .C0(n59), .C1(
        n161), .Y(n1721) );
  XOR2X1TF U1165 ( .A(n1688), .B(n53), .Y(n1140) );
  OAI21X1TF U1166 ( .A0(n2028), .A1(n57), .B0(n1722), .Y(n1688) );
  AOI222XLTF U1167 ( .A0(n49), .A1(n164), .B0(n51), .B1(n161), .C0(n59), .C1(
        n158), .Y(n1722) );
  XOR2X1TF U1168 ( .A(n1689), .B(n53), .Y(n1141) );
  OAI21X1TF U1169 ( .A0(n2029), .A1(n57), .B0(n1723), .Y(n1689) );
  AOI222XLTF U1170 ( .A0(n49), .A1(n161), .B0(n51), .B1(n158), .C0(n59), .C1(
        n155), .Y(n1723) );
  XOR2X1TF U1171 ( .A(n1690), .B(n53), .Y(n1142) );
  OAI21X1TF U1172 ( .A0(n2030), .A1(n56), .B0(n1724), .Y(n1690) );
  AOI222XLTF U1173 ( .A0(n49), .A1(n158), .B0(n51), .B1(n155), .C0(n59), .C1(
        n152), .Y(n1724) );
  XOR2X1TF U1174 ( .A(n1691), .B(n53), .Y(n1143) );
  OAI21X1TF U1175 ( .A0(n2031), .A1(n56), .B0(n1725), .Y(n1691) );
  AOI222XLTF U1176 ( .A0(n49), .A1(n155), .B0(n51), .B1(n152), .C0(n59), .C1(
        n149), .Y(n1725) );
  XOR2X1TF U1177 ( .A(n1692), .B(n53), .Y(n1144) );
  OAI21X1TF U1178 ( .A0(n2032), .A1(n56), .B0(n1726), .Y(n1692) );
  AOI222XLTF U1179 ( .A0(n49), .A1(n152), .B0(n51), .B1(n149), .C0(n59), .C1(
        n146), .Y(n1726) );
  XOR2X1TF U1180 ( .A(n1693), .B(n53), .Y(n1145) );
  OAI21X1TF U1181 ( .A0(n2033), .A1(n56), .B0(n1727), .Y(n1693) );
  AOI222XLTF U1182 ( .A0(n49), .A1(n149), .B0(n51), .B1(n146), .C0(n59), .C1(
        n143), .Y(n1727) );
  XOR2X1TF U1183 ( .A(n1694), .B(n53), .Y(n1146) );
  OAI21X1TF U1184 ( .A0(n2034), .A1(n56), .B0(n1728), .Y(n1694) );
  AOI222XLTF U1185 ( .A0(n49), .A1(n146), .B0(n51), .B1(n143), .C0(n59), .C1(
        n140), .Y(n1728) );
  XOR2X1TF U1186 ( .A(n1695), .B(n53), .Y(n1147) );
  OAI21X1TF U1187 ( .A0(n2035), .A1(n56), .B0(n1729), .Y(n1695) );
  AOI222XLTF U1188 ( .A0(n49), .A1(n143), .B0(n51), .B1(n140), .C0(n59), .C1(
        n137), .Y(n1729) );
  XOR2X1TF U1189 ( .A(n1696), .B(n53), .Y(n1148) );
  OAI21X1TF U1190 ( .A0(n2036), .A1(n56), .B0(n1730), .Y(n1696) );
  AOI222XLTF U1191 ( .A0(n49), .A1(n140), .B0(n51), .B1(n137), .C0(n59), .C1(
        n134), .Y(n1730) );
  XOR2X1TF U1192 ( .A(n1697), .B(n53), .Y(n1149) );
  OAI21X1TF U1193 ( .A0(n2037), .A1(n56), .B0(n1731), .Y(n1697) );
  AOI222XLTF U1194 ( .A0(n49), .A1(n137), .B0(n51), .B1(n134), .C0(n59), .C1(
        n131), .Y(n1731) );
  XOR2X1TF U1195 ( .A(n1698), .B(n53), .Y(n1150) );
  OAI21X1TF U1196 ( .A0(n56), .A1(n2038), .B0(n2294), .Y(n1698) );
  XOR2X1TF U1199 ( .A(n1699), .B(n53), .Y(n1151) );
  OAI21X1TF U1200 ( .A0(n56), .A1(n2039), .B0(n2305), .Y(n1699) );
  INVX2TF U1203 ( .A(n43), .Y(n1152) );
  XOR2X1TF U1204 ( .A(n1734), .B(n43), .Y(n1153) );
  OAI21X1TF U1205 ( .A0(n2006), .A1(n46), .B0(n1768), .Y(n1734) );
  NAND2X1TF U1206 ( .A(n48), .B(n224), .Y(n1768) );
  XOR2X1TF U1207 ( .A(n1735), .B(n43), .Y(n1154) );
  OAI21X1TF U1208 ( .A0(n2007), .A1(n46), .B0(n1769), .Y(n1735) );
  AOI21X1TF U1209 ( .A0(n48), .A1(n221), .B0(n835), .Y(n1769) );
  AND2X2TF U1210 ( .A(n40), .B(n223), .Y(n835) );
  XOR2X1TF U1211 ( .A(n1736), .B(n43), .Y(n1155) );
  OAI21X1TF U1212 ( .A0(n2008), .A1(n46), .B0(n1770), .Y(n1736) );
  AOI222XLTF U1213 ( .A0(n38), .A1(n223), .B0(n40), .B1(n220), .C0(n48), .C1(
        n218), .Y(n1770) );
  XOR2X1TF U1214 ( .A(n1737), .B(n43), .Y(n1156) );
  OAI21X1TF U1215 ( .A0(n2009), .A1(n46), .B0(n1771), .Y(n1737) );
  AOI222XLTF U1216 ( .A0(n38), .A1(n220), .B0(n40), .B1(n217), .C0(n48), .C1(
        n215), .Y(n1771) );
  XOR2X1TF U1217 ( .A(n1738), .B(n43), .Y(n1157) );
  OAI21X1TF U1218 ( .A0(n2010), .A1(n46), .B0(n1772), .Y(n1738) );
  AOI222XLTF U1219 ( .A0(n38), .A1(n217), .B0(n40), .B1(n214), .C0(n48), .C1(
        n212), .Y(n1772) );
  XOR2X1TF U1220 ( .A(n1739), .B(n43), .Y(n1158) );
  OAI21X1TF U1221 ( .A0(n2011), .A1(n46), .B0(n1773), .Y(n1739) );
  AOI222XLTF U1222 ( .A0(n38), .A1(n214), .B0(n40), .B1(n211), .C0(n48), .C1(
        n209), .Y(n1773) );
  XOR2X1TF U1223 ( .A(n1740), .B(n43), .Y(n1159) );
  OAI21X1TF U1224 ( .A0(n2012), .A1(n46), .B0(n1774), .Y(n1740) );
  AOI222XLTF U1225 ( .A0(n38), .A1(n211), .B0(n40), .B1(n208), .C0(n48), .C1(
        n206), .Y(n1774) );
  XOR2X1TF U1226 ( .A(n1741), .B(n43), .Y(n1160) );
  OAI21X1TF U1227 ( .A0(n2013), .A1(n46), .B0(n1775), .Y(n1741) );
  AOI222XLTF U1228 ( .A0(n38), .A1(n208), .B0(n40), .B1(n205), .C0(n48), .C1(
        n203), .Y(n1775) );
  XOR2X1TF U1229 ( .A(n1742), .B(n43), .Y(n1161) );
  OAI21X1TF U1230 ( .A0(n2014), .A1(n46), .B0(n1776), .Y(n1742) );
  AOI222XLTF U1231 ( .A0(n38), .A1(n205), .B0(n40), .B1(n202), .C0(n48), .C1(
        n200), .Y(n1776) );
  XOR2X1TF U1232 ( .A(n1743), .B(n43), .Y(n1162) );
  OAI21X1TF U1233 ( .A0(n2015), .A1(n46), .B0(n1777), .Y(n1743) );
  AOI222XLTF U1234 ( .A0(n38), .A1(n202), .B0(n40), .B1(n199), .C0(n48), .C1(
        n197), .Y(n1777) );
  XOR2X1TF U1235 ( .A(n1744), .B(n42), .Y(n1163) );
  OAI21X1TF U1236 ( .A0(n2016), .A1(n46), .B0(n1778), .Y(n1744) );
  AOI222XLTF U1237 ( .A0(n38), .A1(n199), .B0(n40), .B1(n196), .C0(n48), .C1(
        n194), .Y(n1778) );
  XOR2X1TF U1238 ( .A(n1745), .B(n42), .Y(n1164) );
  OAI21X1TF U1239 ( .A0(n2017), .A1(n46), .B0(n1779), .Y(n1745) );
  AOI222XLTF U1240 ( .A0(n38), .A1(n196), .B0(n40), .B1(n193), .C0(n48), .C1(
        n191), .Y(n1779) );
  XOR2X1TF U1241 ( .A(n1746), .B(n42), .Y(n1165) );
  OAI21X1TF U1242 ( .A0(n2018), .A1(n45), .B0(n1780), .Y(n1746) );
  AOI222XLTF U1243 ( .A0(n38), .A1(n193), .B0(n40), .B1(n190), .C0(n48), .C1(
        n188), .Y(n1780) );
  XOR2X1TF U1244 ( .A(n1747), .B(n42), .Y(n1166) );
  OAI21X1TF U1245 ( .A0(n2019), .A1(n45), .B0(n1781), .Y(n1747) );
  AOI222XLTF U1246 ( .A0(n38), .A1(n190), .B0(n40), .B1(n187), .C0(n48), .C1(
        n185), .Y(n1781) );
  XOR2X1TF U1247 ( .A(n1748), .B(n42), .Y(n1167) );
  OAI21X1TF U1248 ( .A0(n2020), .A1(n45), .B0(n1782), .Y(n1748) );
  AOI222XLTF U1249 ( .A0(n38), .A1(n187), .B0(n40), .B1(n184), .C0(n48), .C1(
        n182), .Y(n1782) );
  XOR2X1TF U1250 ( .A(n1749), .B(n42), .Y(n1168) );
  OAI21X1TF U1251 ( .A0(n2021), .A1(n45), .B0(n1783), .Y(n1749) );
  AOI222XLTF U1252 ( .A0(n38), .A1(n184), .B0(n40), .B1(n181), .C0(n48), .C1(
        n179), .Y(n1783) );
  XOR2X1TF U1253 ( .A(n1750), .B(n42), .Y(n1169) );
  OAI21X1TF U1254 ( .A0(n2022), .A1(n45), .B0(n1784), .Y(n1750) );
  AOI222XLTF U1255 ( .A0(n38), .A1(n181), .B0(n40), .B1(n178), .C0(n47), .C1(
        n176), .Y(n1784) );
  XOR2X1TF U1256 ( .A(n1751), .B(n42), .Y(n1170) );
  OAI21X1TF U1257 ( .A0(n2023), .A1(n45), .B0(n1785), .Y(n1751) );
  AOI222XLTF U1258 ( .A0(n38), .A1(n178), .B0(n39), .B1(n175), .C0(n47), .C1(
        n173), .Y(n1785) );
  XOR2X1TF U1259 ( .A(n1752), .B(n42), .Y(n1171) );
  OAI21X1TF U1260 ( .A0(n2024), .A1(n45), .B0(n1786), .Y(n1752) );
  AOI222XLTF U1261 ( .A0(n37), .A1(n175), .B0(n39), .B1(n172), .C0(n47), .C1(
        n170), .Y(n1786) );
  XOR2X1TF U1262 ( .A(n1753), .B(n42), .Y(n1172) );
  OAI21X1TF U1263 ( .A0(n2025), .A1(n45), .B0(n1787), .Y(n1753) );
  AOI222XLTF U1264 ( .A0(n37), .A1(n172), .B0(n39), .B1(n169), .C0(n47), .C1(
        n167), .Y(n1787) );
  XOR2X1TF U1265 ( .A(n1754), .B(n42), .Y(n1173) );
  OAI21X1TF U1266 ( .A0(n2026), .A1(n45), .B0(n1788), .Y(n1754) );
  AOI222XLTF U1267 ( .A0(n37), .A1(n169), .B0(n39), .B1(n166), .C0(n47), .C1(
        n164), .Y(n1788) );
  XOR2X1TF U1268 ( .A(n1755), .B(n42), .Y(n1174) );
  OAI21X1TF U1269 ( .A0(n2027), .A1(n45), .B0(n1789), .Y(n1755) );
  AOI222XLTF U1270 ( .A0(n37), .A1(n166), .B0(n39), .B1(n163), .C0(n47), .C1(
        n161), .Y(n1789) );
  XOR2X1TF U1271 ( .A(n1756), .B(n41), .Y(n1175) );
  OAI21X1TF U1272 ( .A0(n2028), .A1(n45), .B0(n1790), .Y(n1756) );
  AOI222XLTF U1273 ( .A0(n37), .A1(n163), .B0(n39), .B1(n160), .C0(n47), .C1(
        n158), .Y(n1790) );
  XOR2X1TF U1274 ( .A(n1757), .B(n41), .Y(n1176) );
  OAI21X1TF U1275 ( .A0(n2029), .A1(n45), .B0(n1791), .Y(n1757) );
  AOI222XLTF U1276 ( .A0(n37), .A1(n160), .B0(n39), .B1(n157), .C0(n47), .C1(
        n155), .Y(n1791) );
  XOR2X1TF U1277 ( .A(n1758), .B(n41), .Y(n1177) );
  OAI21X1TF U1278 ( .A0(n2030), .A1(n44), .B0(n1792), .Y(n1758) );
  AOI222XLTF U1279 ( .A0(n37), .A1(n157), .B0(n39), .B1(n154), .C0(n47), .C1(
        n152), .Y(n1792) );
  XOR2X1TF U1280 ( .A(n1759), .B(n41), .Y(n1178) );
  OAI21X1TF U1281 ( .A0(n2031), .A1(n44), .B0(n1793), .Y(n1759) );
  AOI222XLTF U1282 ( .A0(n37), .A1(n154), .B0(n39), .B1(n151), .C0(n47), .C1(
        n149), .Y(n1793) );
  XOR2X1TF U1283 ( .A(n1760), .B(n41), .Y(n1179) );
  OAI21X1TF U1284 ( .A0(n2032), .A1(n44), .B0(n1794), .Y(n1760) );
  AOI222XLTF U1285 ( .A0(n37), .A1(n151), .B0(n39), .B1(n148), .C0(n47), .C1(
        n146), .Y(n1794) );
  XOR2X1TF U1286 ( .A(n1761), .B(n41), .Y(n1180) );
  OAI21X1TF U1287 ( .A0(n2033), .A1(n44), .B0(n1795), .Y(n1761) );
  AOI222XLTF U1288 ( .A0(n37), .A1(n148), .B0(n39), .B1(n145), .C0(n47), .C1(
        n143), .Y(n1795) );
  XOR2X1TF U1289 ( .A(n1762), .B(n41), .Y(n1181) );
  OAI21X1TF U1290 ( .A0(n2034), .A1(n44), .B0(n1796), .Y(n1762) );
  AOI222XLTF U1291 ( .A0(n37), .A1(n145), .B0(n39), .B1(n142), .C0(n47), .C1(
        n140), .Y(n1796) );
  XOR2X1TF U1292 ( .A(n1763), .B(n41), .Y(n1182) );
  OAI21X1TF U1293 ( .A0(n2035), .A1(n44), .B0(n1797), .Y(n1763) );
  AOI222XLTF U1294 ( .A0(n37), .A1(n142), .B0(n39), .B1(n139), .C0(n47), .C1(
        n137), .Y(n1797) );
  XOR2X1TF U1295 ( .A(n1764), .B(n41), .Y(n1183) );
  OAI21X1TF U1296 ( .A0(n2036), .A1(n44), .B0(n1798), .Y(n1764) );
  AOI222XLTF U1297 ( .A0(n37), .A1(n139), .B0(n39), .B1(n136), .C0(n47), .C1(
        n134), .Y(n1798) );
  XOR2X1TF U1298 ( .A(n1765), .B(n41), .Y(n1184) );
  OAI21X1TF U1299 ( .A0(n2037), .A1(n44), .B0(n1799), .Y(n1765) );
  AOI222XLTF U1300 ( .A0(n37), .A1(n136), .B0(n39), .B1(n133), .C0(n47), .C1(
        n131), .Y(n1799) );
  XOR2X1TF U1301 ( .A(n1766), .B(n41), .Y(n1185) );
  OAI21X1TF U1302 ( .A0(n44), .A1(n2038), .B0(n2293), .Y(n1766) );
  XOR2X1TF U1305 ( .A(n1767), .B(n41), .Y(n1186) );
  OAI21X1TF U1306 ( .A0(n44), .A1(n2039), .B0(n2304), .Y(n1767) );
  INVX2TF U1309 ( .A(n31), .Y(n1187) );
  XOR2X1TF U1310 ( .A(n1802), .B(n31), .Y(n1188) );
  OAI21X1TF U1311 ( .A0(n2006), .A1(n34), .B0(n1836), .Y(n1802) );
  NAND2X1TF U1312 ( .A(n36), .B(n223), .Y(n1836) );
  XOR2X1TF U1313 ( .A(n1803), .B(n31), .Y(n1189) );
  OAI21X1TF U1314 ( .A0(n2007), .A1(n34), .B0(n1837), .Y(n1803) );
  AOI21X1TF U1315 ( .A0(n36), .A1(n220), .B0(n838), .Y(n1837) );
  AND2X2TF U1316 ( .A(n28), .B(n223), .Y(n838) );
  XOR2X1TF U1317 ( .A(n1804), .B(n31), .Y(n1190) );
  OAI21X1TF U1318 ( .A0(n2008), .A1(n34), .B0(n1838), .Y(n1804) );
  AOI222XLTF U1319 ( .A0(n26), .A1(n223), .B0(n28), .B1(n220), .C0(n36), .C1(
        n217), .Y(n1838) );
  XOR2X1TF U1320 ( .A(n1805), .B(n31), .Y(n1191) );
  OAI21X1TF U1321 ( .A0(n2009), .A1(n34), .B0(n1839), .Y(n1805) );
  AOI222XLTF U1322 ( .A0(n26), .A1(n220), .B0(n28), .B1(n217), .C0(n36), .C1(
        n214), .Y(n1839) );
  XOR2X1TF U1323 ( .A(n1806), .B(n31), .Y(n1192) );
  OAI21X1TF U1324 ( .A0(n2010), .A1(n34), .B0(n1840), .Y(n1806) );
  AOI222XLTF U1325 ( .A0(n26), .A1(n217), .B0(n28), .B1(n214), .C0(n36), .C1(
        n211), .Y(n1840) );
  XOR2X1TF U1326 ( .A(n1807), .B(n31), .Y(n1193) );
  OAI21X1TF U1327 ( .A0(n2011), .A1(n34), .B0(n1841), .Y(n1807) );
  AOI222XLTF U1328 ( .A0(n26), .A1(n214), .B0(n28), .B1(n211), .C0(n36), .C1(
        n208), .Y(n1841) );
  XOR2X1TF U1329 ( .A(n1808), .B(n31), .Y(n1194) );
  OAI21X1TF U1330 ( .A0(n2012), .A1(n34), .B0(n1842), .Y(n1808) );
  AOI222XLTF U1331 ( .A0(n26), .A1(n211), .B0(n28), .B1(n208), .C0(n36), .C1(
        n205), .Y(n1842) );
  XOR2X1TF U1332 ( .A(n1809), .B(n31), .Y(n1195) );
  OAI21X1TF U1333 ( .A0(n2013), .A1(n34), .B0(n1843), .Y(n1809) );
  AOI222XLTF U1334 ( .A0(n26), .A1(n208), .B0(n28), .B1(n205), .C0(n36), .C1(
        n202), .Y(n1843) );
  XOR2X1TF U1335 ( .A(n1810), .B(n31), .Y(n1196) );
  OAI21X1TF U1336 ( .A0(n2014), .A1(n34), .B0(n1844), .Y(n1810) );
  AOI222XLTF U1337 ( .A0(n26), .A1(n205), .B0(n28), .B1(n202), .C0(n36), .C1(
        n199), .Y(n1844) );
  XOR2X1TF U1338 ( .A(n1811), .B(n31), .Y(n1197) );
  OAI21X1TF U1339 ( .A0(n2015), .A1(n34), .B0(n1845), .Y(n1811) );
  AOI222XLTF U1340 ( .A0(n26), .A1(n202), .B0(n28), .B1(n199), .C0(n36), .C1(
        n196), .Y(n1845) );
  XOR2X1TF U1341 ( .A(n1812), .B(n30), .Y(n1198) );
  OAI21X1TF U1342 ( .A0(n2016), .A1(n34), .B0(n1846), .Y(n1812) );
  AOI222XLTF U1343 ( .A0(n26), .A1(n199), .B0(n28), .B1(n196), .C0(n36), .C1(
        n193), .Y(n1846) );
  XOR2X1TF U1344 ( .A(n1813), .B(n30), .Y(n1199) );
  OAI21X1TF U1345 ( .A0(n2017), .A1(n34), .B0(n1847), .Y(n1813) );
  AOI222XLTF U1346 ( .A0(n26), .A1(n196), .B0(n28), .B1(n193), .C0(n36), .C1(
        n190), .Y(n1847) );
  XOR2X1TF U1347 ( .A(n1814), .B(n30), .Y(n1200) );
  OAI21X1TF U1348 ( .A0(n2018), .A1(n33), .B0(n1848), .Y(n1814) );
  AOI222XLTF U1349 ( .A0(n26), .A1(n193), .B0(n28), .B1(n190), .C0(n36), .C1(
        n187), .Y(n1848) );
  XOR2X1TF U1350 ( .A(n1815), .B(n30), .Y(n1201) );
  OAI21X1TF U1351 ( .A0(n2019), .A1(n33), .B0(n1849), .Y(n1815) );
  AOI222XLTF U1352 ( .A0(n26), .A1(n190), .B0(n28), .B1(n187), .C0(n36), .C1(
        n184), .Y(n1849) );
  XOR2X1TF U1353 ( .A(n1816), .B(n30), .Y(n1202) );
  OAI21X1TF U1354 ( .A0(n2020), .A1(n33), .B0(n1850), .Y(n1816) );
  AOI222XLTF U1355 ( .A0(n26), .A1(n187), .B0(n28), .B1(n184), .C0(n36), .C1(
        n181), .Y(n1850) );
  XOR2X1TF U1356 ( .A(n1817), .B(n30), .Y(n1203) );
  OAI21X1TF U1357 ( .A0(n2021), .A1(n33), .B0(n1851), .Y(n1817) );
  AOI222XLTF U1358 ( .A0(n26), .A1(n184), .B0(n28), .B1(n181), .C0(n36), .C1(
        n178), .Y(n1851) );
  XOR2X1TF U1359 ( .A(n1818), .B(n30), .Y(n1204) );
  OAI21X1TF U1360 ( .A0(n2022), .A1(n33), .B0(n1852), .Y(n1818) );
  AOI222XLTF U1361 ( .A0(n26), .A1(n181), .B0(n28), .B1(n178), .C0(n35), .C1(
        n175), .Y(n1852) );
  XOR2X1TF U1362 ( .A(n1819), .B(n30), .Y(n1205) );
  OAI21X1TF U1363 ( .A0(n2023), .A1(n33), .B0(n1853), .Y(n1819) );
  AOI222XLTF U1364 ( .A0(n26), .A1(n178), .B0(n27), .B1(n175), .C0(n35), .C1(
        n172), .Y(n1853) );
  XOR2X1TF U1365 ( .A(n1820), .B(n30), .Y(n1206) );
  OAI21X1TF U1366 ( .A0(n2024), .A1(n33), .B0(n1854), .Y(n1820) );
  AOI222XLTF U1367 ( .A0(n25), .A1(n175), .B0(n27), .B1(n172), .C0(n35), .C1(
        n169), .Y(n1854) );
  XOR2X1TF U1368 ( .A(n1821), .B(n30), .Y(n1207) );
  OAI21X1TF U1369 ( .A0(n2025), .A1(n33), .B0(n1855), .Y(n1821) );
  AOI222XLTF U1370 ( .A0(n25), .A1(n172), .B0(n27), .B1(n169), .C0(n35), .C1(
        n166), .Y(n1855) );
  XOR2X1TF U1371 ( .A(n1822), .B(n30), .Y(n1208) );
  OAI21X1TF U1372 ( .A0(n2026), .A1(n33), .B0(n1856), .Y(n1822) );
  AOI222XLTF U1373 ( .A0(n25), .A1(n169), .B0(n27), .B1(n166), .C0(n35), .C1(
        n163), .Y(n1856) );
  XOR2X1TF U1374 ( .A(n1823), .B(n30), .Y(n1209) );
  OAI21X1TF U1375 ( .A0(n2027), .A1(n33), .B0(n1857), .Y(n1823) );
  AOI222XLTF U1376 ( .A0(n25), .A1(n166), .B0(n27), .B1(n163), .C0(n35), .C1(
        n160), .Y(n1857) );
  XOR2X1TF U1377 ( .A(n1824), .B(n29), .Y(n1210) );
  OAI21X1TF U1378 ( .A0(n2028), .A1(n33), .B0(n1858), .Y(n1824) );
  AOI222XLTF U1379 ( .A0(n25), .A1(n163), .B0(n27), .B1(n160), .C0(n35), .C1(
        n157), .Y(n1858) );
  XOR2X1TF U1380 ( .A(n1825), .B(n29), .Y(n1211) );
  OAI21X1TF U1381 ( .A0(n2029), .A1(n33), .B0(n1859), .Y(n1825) );
  AOI222XLTF U1382 ( .A0(n25), .A1(n160), .B0(n27), .B1(n157), .C0(n35), .C1(
        n154), .Y(n1859) );
  XOR2X1TF U1383 ( .A(n1826), .B(n29), .Y(n1212) );
  OAI21X1TF U1384 ( .A0(n2030), .A1(n32), .B0(n1860), .Y(n1826) );
  AOI222XLTF U1385 ( .A0(n25), .A1(n157), .B0(n27), .B1(n154), .C0(n35), .C1(
        n151), .Y(n1860) );
  XOR2X1TF U1386 ( .A(n1827), .B(n29), .Y(n1213) );
  OAI21X1TF U1387 ( .A0(n2031), .A1(n32), .B0(n1861), .Y(n1827) );
  AOI222XLTF U1388 ( .A0(n25), .A1(n154), .B0(n27), .B1(n151), .C0(n35), .C1(
        n148), .Y(n1861) );
  XOR2X1TF U1389 ( .A(n1828), .B(n29), .Y(n1214) );
  OAI21X1TF U1390 ( .A0(n2032), .A1(n32), .B0(n1862), .Y(n1828) );
  AOI222XLTF U1391 ( .A0(n25), .A1(n151), .B0(n27), .B1(n148), .C0(n35), .C1(
        n145), .Y(n1862) );
  XOR2X1TF U1392 ( .A(n1829), .B(n29), .Y(n1215) );
  OAI21X1TF U1393 ( .A0(n2033), .A1(n32), .B0(n1863), .Y(n1829) );
  AOI222XLTF U1394 ( .A0(n25), .A1(n148), .B0(n27), .B1(n145), .C0(n35), .C1(
        n142), .Y(n1863) );
  XOR2X1TF U1395 ( .A(n1830), .B(n29), .Y(n1216) );
  OAI21X1TF U1396 ( .A0(n2034), .A1(n32), .B0(n1864), .Y(n1830) );
  AOI222XLTF U1397 ( .A0(n25), .A1(n145), .B0(n27), .B1(n142), .C0(n35), .C1(
        n139), .Y(n1864) );
  XOR2X1TF U1398 ( .A(n1831), .B(n29), .Y(n1217) );
  OAI21X1TF U1399 ( .A0(n2035), .A1(n32), .B0(n1865), .Y(n1831) );
  AOI222XLTF U1400 ( .A0(n25), .A1(n142), .B0(n27), .B1(n139), .C0(n35), .C1(
        n136), .Y(n1865) );
  XOR2X1TF U1401 ( .A(n1832), .B(n29), .Y(n1218) );
  OAI21X1TF U1402 ( .A0(n2036), .A1(n32), .B0(n1866), .Y(n1832) );
  AOI222XLTF U1403 ( .A0(n25), .A1(n139), .B0(n27), .B1(n136), .C0(n35), .C1(
        n133), .Y(n1866) );
  XOR2X1TF U1404 ( .A(n1833), .B(n29), .Y(n1219) );
  OAI21X1TF U1405 ( .A0(n2037), .A1(n32), .B0(n1867), .Y(n1833) );
  AOI222XLTF U1406 ( .A0(n25), .A1(n136), .B0(n27), .B1(n133), .C0(n35), .C1(
        n130), .Y(n1867) );
  XOR2X1TF U1407 ( .A(n1834), .B(n29), .Y(n1220) );
  OAI21X1TF U1408 ( .A0(n32), .A1(n2038), .B0(n2292), .Y(n1834) );
  XOR2X1TF U1411 ( .A(n1835), .B(n29), .Y(n1221) );
  OAI21X1TF U1412 ( .A0(n32), .A1(n2039), .B0(n2303), .Y(n1835) );
  INVX2TF U1415 ( .A(n19), .Y(n1222) );
  XOR2X1TF U1416 ( .A(n1870), .B(n19), .Y(n1223) );
  OAI21X1TF U1417 ( .A0(n2006), .A1(n22), .B0(n1904), .Y(n1870) );
  NAND2X1TF U1418 ( .A(n24), .B(n223), .Y(n1904) );
  XOR2X1TF U1419 ( .A(n1871), .B(n19), .Y(n1224) );
  OAI21X1TF U1420 ( .A0(n2007), .A1(n22), .B0(n1905), .Y(n1871) );
  AOI21X1TF U1421 ( .A0(n24), .A1(n220), .B0(n841), .Y(n1905) );
  AND2X2TF U1422 ( .A(n16), .B(n223), .Y(n841) );
  XOR2X1TF U1423 ( .A(n1872), .B(n19), .Y(n1225) );
  OAI21X1TF U1424 ( .A0(n2008), .A1(n22), .B0(n1906), .Y(n1872) );
  AOI222XLTF U1425 ( .A0(n14), .A1(n223), .B0(n16), .B1(n220), .C0(n24), .C1(
        n217), .Y(n1906) );
  XOR2X1TF U1426 ( .A(n1873), .B(n19), .Y(n1226) );
  OAI21X1TF U1427 ( .A0(n2009), .A1(n22), .B0(n1907), .Y(n1873) );
  AOI222XLTF U1428 ( .A0(n14), .A1(n220), .B0(n16), .B1(n217), .C0(n24), .C1(
        n214), .Y(n1907) );
  XOR2X1TF U1429 ( .A(n1874), .B(n19), .Y(n1227) );
  OAI21X1TF U1430 ( .A0(n2010), .A1(n22), .B0(n1908), .Y(n1874) );
  AOI222XLTF U1431 ( .A0(n14), .A1(n217), .B0(n16), .B1(n214), .C0(n24), .C1(
        n211), .Y(n1908) );
  XOR2X1TF U1432 ( .A(n1875), .B(n19), .Y(n1228) );
  OAI21X1TF U1433 ( .A0(n2011), .A1(n22), .B0(n1909), .Y(n1875) );
  AOI222XLTF U1434 ( .A0(n14), .A1(n214), .B0(n16), .B1(n211), .C0(n24), .C1(
        n208), .Y(n1909) );
  XOR2X1TF U1435 ( .A(n1876), .B(n19), .Y(n1229) );
  OAI21X1TF U1436 ( .A0(n2012), .A1(n22), .B0(n1910), .Y(n1876) );
  AOI222XLTF U1437 ( .A0(n14), .A1(n211), .B0(n16), .B1(n208), .C0(n24), .C1(
        n205), .Y(n1910) );
  XOR2X1TF U1438 ( .A(n1877), .B(n19), .Y(n1230) );
  OAI21X1TF U1439 ( .A0(n2013), .A1(n22), .B0(n1911), .Y(n1877) );
  AOI222XLTF U1440 ( .A0(n14), .A1(n208), .B0(n16), .B1(n205), .C0(n24), .C1(
        n202), .Y(n1911) );
  XOR2X1TF U1441 ( .A(n1878), .B(n19), .Y(n1231) );
  OAI21X1TF U1442 ( .A0(n2014), .A1(n22), .B0(n1912), .Y(n1878) );
  AOI222XLTF U1443 ( .A0(n14), .A1(n205), .B0(n16), .B1(n202), .C0(n24), .C1(
        n199), .Y(n1912) );
  XOR2X1TF U1444 ( .A(n1879), .B(n19), .Y(n1232) );
  OAI21X1TF U1445 ( .A0(n2015), .A1(n22), .B0(n1913), .Y(n1879) );
  AOI222XLTF U1446 ( .A0(n14), .A1(n202), .B0(n16), .B1(n199), .C0(n24), .C1(
        n196), .Y(n1913) );
  XOR2X1TF U1447 ( .A(n1880), .B(n18), .Y(n1233) );
  OAI21X1TF U1448 ( .A0(n2016), .A1(n22), .B0(n1914), .Y(n1880) );
  AOI222XLTF U1449 ( .A0(n14), .A1(n199), .B0(n16), .B1(n196), .C0(n24), .C1(
        n193), .Y(n1914) );
  XOR2X1TF U1450 ( .A(n1881), .B(n18), .Y(n1234) );
  OAI21X1TF U1451 ( .A0(n2017), .A1(n22), .B0(n1915), .Y(n1881) );
  AOI222XLTF U1452 ( .A0(n14), .A1(n196), .B0(n16), .B1(n193), .C0(n24), .C1(
        n190), .Y(n1915) );
  XOR2X1TF U1453 ( .A(n1882), .B(n18), .Y(n1235) );
  OAI21X1TF U1454 ( .A0(n2018), .A1(n21), .B0(n1916), .Y(n1882) );
  AOI222XLTF U1455 ( .A0(n14), .A1(n193), .B0(n16), .B1(n190), .C0(n24), .C1(
        n187), .Y(n1916) );
  XOR2X1TF U1456 ( .A(n1883), .B(n18), .Y(n1236) );
  OAI21X1TF U1457 ( .A0(n2019), .A1(n21), .B0(n1917), .Y(n1883) );
  AOI222XLTF U1458 ( .A0(n14), .A1(n190), .B0(n16), .B1(n187), .C0(n24), .C1(
        n184), .Y(n1917) );
  XOR2X1TF U1459 ( .A(n1884), .B(n18), .Y(n1237) );
  OAI21X1TF U1460 ( .A0(n2020), .A1(n21), .B0(n1918), .Y(n1884) );
  AOI222XLTF U1461 ( .A0(n14), .A1(n187), .B0(n16), .B1(n184), .C0(n24), .C1(
        n181), .Y(n1918) );
  XOR2X1TF U1462 ( .A(n1885), .B(n18), .Y(n1238) );
  OAI21X1TF U1463 ( .A0(n2021), .A1(n21), .B0(n1919), .Y(n1885) );
  AOI222XLTF U1464 ( .A0(n14), .A1(n184), .B0(n16), .B1(n181), .C0(n24), .C1(
        n178), .Y(n1919) );
  XOR2X1TF U1465 ( .A(n1886), .B(n18), .Y(n1239) );
  OAI21X1TF U1466 ( .A0(n2022), .A1(n21), .B0(n1920), .Y(n1886) );
  AOI222XLTF U1467 ( .A0(n14), .A1(n181), .B0(n16), .B1(n178), .C0(n23), .C1(
        n175), .Y(n1920) );
  XOR2X1TF U1468 ( .A(n1887), .B(n18), .Y(n1240) );
  OAI21X1TF U1469 ( .A0(n2023), .A1(n21), .B0(n1921), .Y(n1887) );
  AOI222XLTF U1470 ( .A0(n14), .A1(n178), .B0(n15), .B1(n175), .C0(n23), .C1(
        n172), .Y(n1921) );
  XOR2X1TF U1471 ( .A(n1888), .B(n18), .Y(n1241) );
  OAI21X1TF U1472 ( .A0(n2024), .A1(n21), .B0(n1922), .Y(n1888) );
  AOI222XLTF U1473 ( .A0(n13), .A1(n175), .B0(n15), .B1(n172), .C0(n23), .C1(
        n169), .Y(n1922) );
  XOR2X1TF U1474 ( .A(n1889), .B(n18), .Y(n1242) );
  OAI21X1TF U1475 ( .A0(n2025), .A1(n21), .B0(n1923), .Y(n1889) );
  AOI222XLTF U1476 ( .A0(n13), .A1(n172), .B0(n15), .B1(n169), .C0(n23), .C1(
        n166), .Y(n1923) );
  XOR2X1TF U1477 ( .A(n1890), .B(n18), .Y(n1243) );
  OAI21X1TF U1478 ( .A0(n2026), .A1(n21), .B0(n1924), .Y(n1890) );
  AOI222XLTF U1479 ( .A0(n13), .A1(n169), .B0(n15), .B1(n166), .C0(n23), .C1(
        n163), .Y(n1924) );
  XOR2X1TF U1480 ( .A(n1891), .B(n18), .Y(n1244) );
  OAI21X1TF U1481 ( .A0(n2027), .A1(n21), .B0(n1925), .Y(n1891) );
  AOI222XLTF U1482 ( .A0(n13), .A1(n166), .B0(n15), .B1(n163), .C0(n23), .C1(
        n160), .Y(n1925) );
  XOR2X1TF U1483 ( .A(n1892), .B(n17), .Y(n1245) );
  OAI21X1TF U1484 ( .A0(n2028), .A1(n21), .B0(n1926), .Y(n1892) );
  AOI222XLTF U1485 ( .A0(n13), .A1(n163), .B0(n15), .B1(n160), .C0(n23), .C1(
        n157), .Y(n1926) );
  XOR2X1TF U1486 ( .A(n1893), .B(n17), .Y(n1246) );
  OAI21X1TF U1487 ( .A0(n2029), .A1(n21), .B0(n1927), .Y(n1893) );
  AOI222XLTF U1488 ( .A0(n13), .A1(n160), .B0(n15), .B1(n157), .C0(n23), .C1(
        n154), .Y(n1927) );
  XOR2X1TF U1489 ( .A(n1894), .B(n17), .Y(n1247) );
  OAI21X1TF U1490 ( .A0(n2030), .A1(n20), .B0(n1928), .Y(n1894) );
  AOI222XLTF U1491 ( .A0(n13), .A1(n157), .B0(n15), .B1(n154), .C0(n23), .C1(
        n151), .Y(n1928) );
  XOR2X1TF U1492 ( .A(n1895), .B(n17), .Y(n1248) );
  OAI21X1TF U1493 ( .A0(n2031), .A1(n20), .B0(n1929), .Y(n1895) );
  AOI222XLTF U1494 ( .A0(n13), .A1(n154), .B0(n15), .B1(n151), .C0(n23), .C1(
        n148), .Y(n1929) );
  XOR2X1TF U1495 ( .A(n1896), .B(n17), .Y(n1249) );
  OAI21X1TF U1496 ( .A0(n2032), .A1(n20), .B0(n1930), .Y(n1896) );
  AOI222XLTF U1497 ( .A0(n13), .A1(n151), .B0(n15), .B1(n148), .C0(n23), .C1(
        n145), .Y(n1930) );
  XOR2X1TF U1498 ( .A(n1897), .B(n17), .Y(n1250) );
  OAI21X1TF U1499 ( .A0(n2033), .A1(n20), .B0(n1931), .Y(n1897) );
  AOI222XLTF U1500 ( .A0(n13), .A1(n148), .B0(n15), .B1(n145), .C0(n23), .C1(
        n142), .Y(n1931) );
  XOR2X1TF U1501 ( .A(n1898), .B(n17), .Y(n1251) );
  OAI21X1TF U1502 ( .A0(n2034), .A1(n20), .B0(n1932), .Y(n1898) );
  AOI222XLTF U1503 ( .A0(n13), .A1(n145), .B0(n15), .B1(n142), .C0(n23), .C1(
        n139), .Y(n1932) );
  XOR2X1TF U1504 ( .A(n1899), .B(n17), .Y(n1252) );
  OAI21X1TF U1505 ( .A0(n2035), .A1(n20), .B0(n1933), .Y(n1899) );
  AOI222XLTF U1506 ( .A0(n13), .A1(n142), .B0(n15), .B1(n139), .C0(n23), .C1(
        n136), .Y(n1933) );
  XOR2X1TF U1507 ( .A(n1900), .B(n17), .Y(n1253) );
  OAI21X1TF U1508 ( .A0(n2036), .A1(n20), .B0(n1934), .Y(n1900) );
  AOI222XLTF U1509 ( .A0(n13), .A1(n139), .B0(n15), .B1(n136), .C0(n23), .C1(
        n133), .Y(n1934) );
  XOR2X1TF U1510 ( .A(n1901), .B(n17), .Y(n1254) );
  OAI21X1TF U1511 ( .A0(n2037), .A1(n20), .B0(n1935), .Y(n1901) );
  AOI222XLTF U1512 ( .A0(n13), .A1(n136), .B0(n15), .B1(n133), .C0(n23), .C1(
        n130), .Y(n1935) );
  XOR2X1TF U1513 ( .A(n1902), .B(n17), .Y(n1255) );
  OAI21X1TF U1514 ( .A0(n20), .A1(n2038), .B0(n2291), .Y(n1902) );
  XOR2X1TF U1517 ( .A(n1903), .B(n17), .Y(n1256) );
  OAI21X1TF U1518 ( .A0(n20), .A1(n2039), .B0(n2302), .Y(n1903) );
  INVX2TF U1521 ( .A(n7), .Y(n1257) );
  XOR2X1TF U1522 ( .A(n1938), .B(n7), .Y(n1258) );
  OAI21X1TF U1523 ( .A0(n2006), .A1(n10), .B0(n1972), .Y(n1938) );
  NAND2X1TF U1524 ( .A(n12), .B(n223), .Y(n1972) );
  XOR2X1TF U1525 ( .A(n1939), .B(n7), .Y(n1259) );
  OAI21X1TF U1526 ( .A0(n2007), .A1(n10), .B0(n1973), .Y(n1939) );
  AOI21X1TF U1527 ( .A0(n12), .A1(n220), .B0(n844), .Y(n1973) );
  AND2X2TF U1528 ( .A(n4), .B(n223), .Y(n844) );
  XOR2X1TF U1529 ( .A(n1940), .B(n7), .Y(n1260) );
  OAI21X1TF U1530 ( .A0(n2008), .A1(n10), .B0(n1974), .Y(n1940) );
  AOI222XLTF U1531 ( .A0(n2), .A1(n223), .B0(n4), .B1(n220), .C0(n12), .C1(
        n217), .Y(n1974) );
  XOR2X1TF U1532 ( .A(n1941), .B(n7), .Y(n1261) );
  OAI21X1TF U1533 ( .A0(n2009), .A1(n10), .B0(n1975), .Y(n1941) );
  AOI222XLTF U1534 ( .A0(n2), .A1(n220), .B0(n4), .B1(n217), .C0(n12), .C1(
        n214), .Y(n1975) );
  XOR2X1TF U1535 ( .A(n1942), .B(n7), .Y(n1262) );
  OAI21X1TF U1536 ( .A0(n2010), .A1(n10), .B0(n1976), .Y(n1942) );
  AOI222XLTF U1537 ( .A0(n2), .A1(n217), .B0(n4), .B1(n214), .C0(n12), .C1(
        n211), .Y(n1976) );
  XOR2X1TF U1538 ( .A(n1943), .B(n7), .Y(n1263) );
  OAI21X1TF U1539 ( .A0(n2011), .A1(n10), .B0(n1977), .Y(n1943) );
  AOI222XLTF U1540 ( .A0(n2), .A1(n214), .B0(n4), .B1(n211), .C0(n12), .C1(
        n208), .Y(n1977) );
  XOR2X1TF U1541 ( .A(n1944), .B(n7), .Y(n1264) );
  OAI21X1TF U1542 ( .A0(n2012), .A1(n10), .B0(n1978), .Y(n1944) );
  AOI222XLTF U1543 ( .A0(n2), .A1(n211), .B0(n4), .B1(n208), .C0(n12), .C1(
        n205), .Y(n1978) );
  XOR2X1TF U1544 ( .A(n1945), .B(n7), .Y(n1265) );
  OAI21X1TF U1545 ( .A0(n2013), .A1(n10), .B0(n1979), .Y(n1945) );
  AOI222XLTF U1546 ( .A0(n2), .A1(n208), .B0(n4), .B1(n205), .C0(n12), .C1(
        n202), .Y(n1979) );
  XOR2X1TF U1547 ( .A(n1946), .B(n6), .Y(n1266) );
  OAI21X1TF U1548 ( .A0(n2014), .A1(n10), .B0(n1980), .Y(n1946) );
  AOI222XLTF U1549 ( .A0(n2), .A1(n205), .B0(n4), .B1(n202), .C0(n12), .C1(
        n199), .Y(n1980) );
  XOR2X1TF U1550 ( .A(n1947), .B(n6), .Y(n1267) );
  OAI21X1TF U1551 ( .A0(n2015), .A1(n10), .B0(n1981), .Y(n1947) );
  AOI222XLTF U1552 ( .A0(n2), .A1(n202), .B0(n4), .B1(n199), .C0(n12), .C1(
        n196), .Y(n1981) );
  XOR2X1TF U1553 ( .A(n1948), .B(n6), .Y(n1268) );
  OAI21X1TF U1554 ( .A0(n2016), .A1(n10), .B0(n1982), .Y(n1948) );
  AOI222XLTF U1555 ( .A0(n2), .A1(n199), .B0(n4), .B1(n196), .C0(n12), .C1(
        n193), .Y(n1982) );
  XOR2X1TF U1556 ( .A(n1949), .B(n6), .Y(n1269) );
  OAI21X1TF U1557 ( .A0(n2017), .A1(n10), .B0(n1983), .Y(n1949) );
  AOI222XLTF U1558 ( .A0(n2), .A1(n196), .B0(n4), .B1(n193), .C0(n12), .C1(
        n190), .Y(n1983) );
  XOR2X1TF U1559 ( .A(n1950), .B(n6), .Y(n1270) );
  OAI21X1TF U1560 ( .A0(n2018), .A1(n9), .B0(n1984), .Y(n1950) );
  AOI222XLTF U1561 ( .A0(n2), .A1(n193), .B0(n4), .B1(n190), .C0(n12), .C1(
        n187), .Y(n1984) );
  XOR2X1TF U1562 ( .A(n1951), .B(n6), .Y(n1271) );
  OAI21X1TF U1563 ( .A0(n2019), .A1(n9), .B0(n1985), .Y(n1951) );
  AOI222XLTF U1564 ( .A0(n2), .A1(n190), .B0(n4), .B1(n187), .C0(n12), .C1(
        n184), .Y(n1985) );
  XOR2X1TF U1565 ( .A(n1952), .B(n6), .Y(n1272) );
  OAI21X1TF U1566 ( .A0(n2020), .A1(n9), .B0(n1986), .Y(n1952) );
  AOI222XLTF U1567 ( .A0(n2), .A1(n187), .B0(n4), .B1(n184), .C0(n12), .C1(
        n181), .Y(n1986) );
  XOR2X1TF U1568 ( .A(n1953), .B(n6), .Y(n1273) );
  OAI21X1TF U1569 ( .A0(n2021), .A1(n9), .B0(n1987), .Y(n1953) );
  AOI222XLTF U1570 ( .A0(n2), .A1(n184), .B0(n4), .B1(n181), .C0(n12), .C1(
        n178), .Y(n1987) );
  XOR2X1TF U1571 ( .A(n1954), .B(n6), .Y(n1274) );
  OAI21X1TF U1572 ( .A0(n2022), .A1(n9), .B0(n1988), .Y(n1954) );
  AOI222XLTF U1573 ( .A0(n2), .A1(n181), .B0(n4), .B1(n178), .C0(n11), .C1(
        n175), .Y(n1988) );
  XOR2X1TF U1574 ( .A(n1955), .B(n6), .Y(n1275) );
  OAI21X1TF U1575 ( .A0(n2023), .A1(n9), .B0(n1989), .Y(n1955) );
  AOI222XLTF U1576 ( .A0(n2), .A1(n178), .B0(n3), .B1(n175), .C0(n11), .C1(
        n172), .Y(n1989) );
  XOR2X1TF U1577 ( .A(n1956), .B(n6), .Y(n1276) );
  OAI21X1TF U1578 ( .A0(n2024), .A1(n9), .B0(n1990), .Y(n1956) );
  AOI222XLTF U1579 ( .A0(n1), .A1(n175), .B0(n3), .B1(n172), .C0(n11), .C1(
        n169), .Y(n1990) );
  XOR2X1TF U1580 ( .A(n1957), .B(n6), .Y(n1277) );
  OAI21X1TF U1581 ( .A0(n2025), .A1(n9), .B0(n1991), .Y(n1957) );
  AOI222XLTF U1582 ( .A0(n1), .A1(n172), .B0(n3), .B1(n169), .C0(n11), .C1(
        n166), .Y(n1991) );
  XOR2X1TF U1583 ( .A(n1958), .B(n6), .Y(n1278) );
  OAI21X1TF U1584 ( .A0(n2026), .A1(n9), .B0(n1992), .Y(n1958) );
  AOI222XLTF U1585 ( .A0(n1), .A1(n169), .B0(n3), .B1(n166), .C0(n11), .C1(
        n163), .Y(n1992) );
  XOR2X1TF U1586 ( .A(n1959), .B(n5), .Y(n1279) );
  OAI21X1TF U1587 ( .A0(n2027), .A1(n9), .B0(n1993), .Y(n1959) );
  AOI222XLTF U1588 ( .A0(n1), .A1(n166), .B0(n3), .B1(n163), .C0(n11), .C1(
        n160), .Y(n1993) );
  XOR2X1TF U1589 ( .A(n1960), .B(n5), .Y(n1280) );
  OAI21X1TF U1590 ( .A0(n2028), .A1(n9), .B0(n1994), .Y(n1960) );
  AOI222XLTF U1591 ( .A0(n1), .A1(n163), .B0(n3), .B1(n160), .C0(n11), .C1(
        n157), .Y(n1994) );
  XOR2X1TF U1592 ( .A(n1961), .B(n5), .Y(n1281) );
  OAI21X1TF U1593 ( .A0(n2029), .A1(n9), .B0(n1995), .Y(n1961) );
  AOI222XLTF U1594 ( .A0(n1), .A1(n160), .B0(n3), .B1(n157), .C0(n11), .C1(
        n154), .Y(n1995) );
  XOR2X1TF U1595 ( .A(n1962), .B(n5), .Y(n1282) );
  OAI21X1TF U1596 ( .A0(n2030), .A1(n8), .B0(n1996), .Y(n1962) );
  AOI222XLTF U1597 ( .A0(n1), .A1(n157), .B0(n3), .B1(n154), .C0(n11), .C1(
        n151), .Y(n1996) );
  XOR2X1TF U1598 ( .A(n1963), .B(n5), .Y(n1283) );
  OAI21X1TF U1599 ( .A0(n2031), .A1(n8), .B0(n1997), .Y(n1963) );
  AOI222XLTF U1600 ( .A0(n1), .A1(n154), .B0(n3), .B1(n151), .C0(n11), .C1(
        n148), .Y(n1997) );
  XOR2X1TF U1601 ( .A(n1964), .B(n5), .Y(n1284) );
  OAI21X1TF U1602 ( .A0(n2032), .A1(n8), .B0(n1998), .Y(n1964) );
  AOI222XLTF U1603 ( .A0(n1), .A1(n151), .B0(n3), .B1(n148), .C0(n11), .C1(
        n145), .Y(n1998) );
  XOR2X1TF U1604 ( .A(n1965), .B(n5), .Y(n1285) );
  OAI21X1TF U1605 ( .A0(n2033), .A1(n8), .B0(n1999), .Y(n1965) );
  AOI222XLTF U1606 ( .A0(n1), .A1(n148), .B0(n3), .B1(n145), .C0(n11), .C1(
        n142), .Y(n1999) );
  XOR2X1TF U1607 ( .A(n1966), .B(n5), .Y(n1286) );
  OAI21X1TF U1608 ( .A0(n2034), .A1(n8), .B0(n2000), .Y(n1966) );
  AOI222XLTF U1609 ( .A0(n1), .A1(n145), .B0(n3), .B1(n142), .C0(n11), .C1(
        n139), .Y(n2000) );
  XOR2X1TF U1610 ( .A(n1967), .B(n5), .Y(n1287) );
  OAI21X1TF U1611 ( .A0(n2035), .A1(n8), .B0(n2001), .Y(n1967) );
  AOI222XLTF U1612 ( .A0(n1), .A1(n142), .B0(n3), .B1(n139), .C0(n11), .C1(
        n136), .Y(n2001) );
  XOR2X1TF U1613 ( .A(n1968), .B(n5), .Y(n1288) );
  OAI21X1TF U1614 ( .A0(n2036), .A1(n8), .B0(n2002), .Y(n1968) );
  AOI222XLTF U1615 ( .A0(n1), .A1(n139), .B0(n3), .B1(n136), .C0(n11), .C1(
        n133), .Y(n2002) );
  XOR2X1TF U1616 ( .A(n1969), .B(n5), .Y(n1289) );
  OAI21X1TF U1617 ( .A0(n2037), .A1(n8), .B0(n2003), .Y(n1969) );
  AOI222XLTF U1618 ( .A0(n1), .A1(n136), .B0(n3), .B1(n133), .C0(n11), .C1(
        n130), .Y(n2003) );
  XOR2X1TF U1619 ( .A(n1970), .B(n5), .Y(n1290) );
  OAI21X1TF U1620 ( .A0(n2038), .A1(n8), .B0(n2290), .Y(n1970) );
  XOR2X1TF U1623 ( .A(n1971), .B(n5), .Y(n1291) );
  OAI21X1TF U1624 ( .A0(n8), .A1(n2039), .B0(n2301), .Y(n1971) );
  AND3X2TF U1703 ( .A(n2072), .B(n2083), .C(a[31]), .Y(n2105) );
  NAND2BX1TF U1704 ( .AN(n2072), .B(a[31]), .Y(n2116) );
  NOR2BX1TF U1705 ( .AN(n2072), .B(n2083), .Y(n2127) );
  NOR2X1TF U1706 ( .A(n2072), .B(a[31]), .Y(n2138) );
  XNOR2X1TF U1707 ( .A(a[30]), .B(a[31]), .Y(n2083) );
  XNOR2X1TF U1708 ( .A(a[29]), .B(a[30]), .Y(n2072) );
  AND3X2TF U1709 ( .A(n2073), .B(n2084), .C(n2095), .Y(n2106) );
  NAND2BX1TF U1710 ( .AN(n2073), .B(n2095), .Y(n2117) );
  NOR2BX1TF U1711 ( .AN(n2073), .B(n2084), .Y(n2128) );
  NOR2X1TF U1712 ( .A(n2073), .B(n2095), .Y(n2139) );
  XNOR2X1TF U1713 ( .A(a[27]), .B(a[28]), .Y(n2084) );
  XNOR2X1TF U1714 ( .A(a[26]), .B(a[27]), .Y(n2073) );
  XOR2X1TF U1715 ( .A(a[28]), .B(a[29]), .Y(n2095) );
  AND3X2TF U1716 ( .A(n2074), .B(n2085), .C(n2096), .Y(n2107) );
  NAND2BX1TF U1717 ( .AN(n2074), .B(n2096), .Y(n2118) );
  NOR2BX1TF U1718 ( .AN(n2074), .B(n2085), .Y(n2129) );
  NOR2X1TF U1719 ( .A(n2074), .B(n2096), .Y(n2140) );
  XNOR2X1TF U1720 ( .A(a[24]), .B(a[25]), .Y(n2085) );
  XNOR2X1TF U1721 ( .A(a[23]), .B(a[24]), .Y(n2074) );
  XOR2X1TF U1722 ( .A(a[25]), .B(a[26]), .Y(n2096) );
  AND3X2TF U1723 ( .A(n2075), .B(n2086), .C(n2097), .Y(n2108) );
  NAND2BX1TF U1724 ( .AN(n2075), .B(n2097), .Y(n2119) );
  NOR2BX1TF U1725 ( .AN(n2075), .B(n2086), .Y(n2130) );
  NOR2X1TF U1726 ( .A(n2075), .B(n2097), .Y(n2141) );
  XNOR2X1TF U1727 ( .A(a[21]), .B(a[22]), .Y(n2086) );
  XNOR2X1TF U1728 ( .A(a[20]), .B(a[21]), .Y(n2075) );
  XOR2X1TF U1729 ( .A(a[22]), .B(a[23]), .Y(n2097) );
  AND3X2TF U1730 ( .A(n2076), .B(n2087), .C(n2098), .Y(n2109) );
  NAND2BX1TF U1731 ( .AN(n2076), .B(n2098), .Y(n2120) );
  NOR2BX1TF U1732 ( .AN(n2076), .B(n2087), .Y(n2131) );
  NOR2X1TF U1733 ( .A(n2076), .B(n2098), .Y(n2142) );
  XNOR2X1TF U1734 ( .A(a[18]), .B(a[19]), .Y(n2087) );
  XNOR2X1TF U1735 ( .A(a[17]), .B(a[18]), .Y(n2076) );
  XOR2X1TF U1736 ( .A(a[19]), .B(a[20]), .Y(n2098) );
  AND3X2TF U1737 ( .A(n2077), .B(n2088), .C(n2099), .Y(n2110) );
  NAND2BX1TF U1738 ( .AN(n2077), .B(n2099), .Y(n2121) );
  NOR2BX1TF U1739 ( .AN(n2077), .B(n2088), .Y(n2132) );
  NOR2X1TF U1740 ( .A(n2077), .B(n2099), .Y(n2143) );
  XNOR2X1TF U1741 ( .A(a[15]), .B(a[16]), .Y(n2088) );
  XNOR2X1TF U1742 ( .A(a[14]), .B(a[15]), .Y(n2077) );
  XOR2X1TF U1743 ( .A(a[16]), .B(a[17]), .Y(n2099) );
  AND3X2TF U1744 ( .A(n2078), .B(n2089), .C(n2100), .Y(n2111) );
  NAND2BX1TF U1745 ( .AN(n2078), .B(n2100), .Y(n2122) );
  NOR2BX1TF U1746 ( .AN(n2078), .B(n2089), .Y(n2133) );
  NOR2X1TF U1747 ( .A(n2078), .B(n2100), .Y(n2144) );
  XNOR2X1TF U1748 ( .A(a[12]), .B(a[13]), .Y(n2089) );
  XNOR2X1TF U1749 ( .A(a[11]), .B(a[12]), .Y(n2078) );
  XOR2X1TF U1750 ( .A(a[13]), .B(a[14]), .Y(n2100) );
  AND3X2TF U1751 ( .A(n2079), .B(n2090), .C(n2101), .Y(n2112) );
  NAND2BX1TF U1752 ( .AN(n2079), .B(n2101), .Y(n2123) );
  NOR2BX1TF U1753 ( .AN(n2079), .B(n2090), .Y(n2134) );
  NOR2X1TF U1754 ( .A(n2079), .B(n2101), .Y(n2145) );
  XNOR2X1TF U1755 ( .A(a[9]), .B(a[10]), .Y(n2090) );
  XNOR2X1TF U1756 ( .A(a[8]), .B(a[9]), .Y(n2079) );
  XOR2X1TF U1757 ( .A(a[10]), .B(a[11]), .Y(n2101) );
  AND3X2TF U1758 ( .A(n2080), .B(n2091), .C(n2102), .Y(n2113) );
  NAND2BX1TF U1759 ( .AN(n2080), .B(n2102), .Y(n2124) );
  NOR2BX1TF U1760 ( .AN(n2080), .B(n2091), .Y(n2135) );
  NOR2X1TF U1761 ( .A(n2080), .B(n2102), .Y(n2146) );
  XNOR2X1TF U1762 ( .A(a[6]), .B(a[7]), .Y(n2091) );
  XNOR2X1TF U1763 ( .A(a[5]), .B(a[6]), .Y(n2080) );
  XOR2X1TF U1764 ( .A(a[7]), .B(a[8]), .Y(n2102) );
  AND3X2TF U1765 ( .A(n2081), .B(n2092), .C(n2103), .Y(n2114) );
  NAND2BX1TF U1766 ( .AN(n2081), .B(n2103), .Y(n2125) );
  NOR2BX1TF U1767 ( .AN(n2081), .B(n2092), .Y(n2136) );
  NOR2X1TF U1768 ( .A(n2081), .B(n2103), .Y(n2147) );
  XNOR2X1TF U1769 ( .A(a[3]), .B(a[4]), .Y(n2092) );
  XNOR2X1TF U1770 ( .A(a[2]), .B(a[3]), .Y(n2081) );
  XOR2X1TF U1771 ( .A(a[4]), .B(a[5]), .Y(n2103) );
  AND3X2TF U1772 ( .A(n2093), .B(n2104), .C(n2082), .Y(n2115) );
  NAND2BX1TF U1773 ( .AN(n2082), .B(n2104), .Y(n2126) );
  NOR2BX1TF U1774 ( .AN(n2082), .B(n2093), .Y(n2137) );
  NOR2X1TF U1775 ( .A(n2104), .B(n2082), .Y(n2148) );
  XNOR2X1TF U1776 ( .A(a[0]), .B(a[1]), .Y(n2093) );
  INVX2TF U1777 ( .A(a[0]), .Y(n2082) );
  XOR2X1TF U1778 ( .A(a[1]), .B(a[2]), .Y(n2104) );
  ADDHXLTF U1779 ( .A(b[31]), .B(n847), .CO(n878), .S(n879) );
  CMPR32X2TF U1780 ( .A(b[30]), .B(b[31]), .C(n848), .CO(n847), .S(n880) );
  CMPR32X2TF U1781 ( .A(b[29]), .B(b[30]), .C(n849), .CO(n848), .S(n881) );
  CMPR32X2TF U1782 ( .A(b[28]), .B(b[29]), .C(n850), .CO(n849), .S(n882) );
  CMPR32X2TF U1783 ( .A(b[27]), .B(b[28]), .C(n851), .CO(n850), .S(n883) );
  CMPR32X2TF U1784 ( .A(b[26]), .B(b[27]), .C(n852), .CO(n851), .S(n884) );
  CMPR32X2TF U1785 ( .A(b[25]), .B(b[26]), .C(n853), .CO(n852), .S(n885) );
  CMPR32X2TF U1786 ( .A(b[24]), .B(b[25]), .C(n854), .CO(n853), .S(n886) );
  CMPR32X2TF U1787 ( .A(b[23]), .B(b[24]), .C(n855), .CO(n854), .S(n887) );
  CMPR32X2TF U1788 ( .A(b[22]), .B(b[23]), .C(n856), .CO(n855), .S(n888) );
  CMPR32X2TF U1789 ( .A(b[21]), .B(b[22]), .C(n857), .CO(n856), .S(n889) );
  CMPR32X2TF U1790 ( .A(b[20]), .B(b[21]), .C(n858), .CO(n857), .S(n890) );
  CMPR32X2TF U1791 ( .A(b[19]), .B(b[20]), .C(n859), .CO(n858), .S(n891) );
  CMPR32X2TF U1792 ( .A(b[18]), .B(b[19]), .C(n860), .CO(n859), .S(n892) );
  CMPR32X2TF U1793 ( .A(b[17]), .B(b[18]), .C(n861), .CO(n860), .S(n893) );
  CMPR32X2TF U1794 ( .A(b[16]), .B(b[17]), .C(n862), .CO(n861), .S(n894) );
  CMPR32X2TF U1795 ( .A(b[15]), .B(b[16]), .C(n863), .CO(n862), .S(n895) );
  CMPR32X2TF U1796 ( .A(b[14]), .B(b[15]), .C(n864), .CO(n863), .S(n896) );
  CMPR32X2TF U1797 ( .A(b[13]), .B(b[14]), .C(n865), .CO(n864), .S(n897) );
  CMPR32X2TF U1798 ( .A(b[12]), .B(b[13]), .C(n866), .CO(n865), .S(n898) );
  CMPR32X2TF U1799 ( .A(b[11]), .B(b[12]), .C(n867), .CO(n866), .S(n899) );
  CMPR32X2TF U1800 ( .A(b[10]), .B(b[11]), .C(n868), .CO(n867), .S(n900) );
  CMPR32X2TF U1801 ( .A(b[9]), .B(b[10]), .C(n869), .CO(n868), .S(n901) );
  CMPR32X2TF U1802 ( .A(b[8]), .B(b[9]), .C(n870), .CO(n869), .S(n902) );
  CMPR32X2TF U1803 ( .A(b[7]), .B(b[8]), .C(n871), .CO(n870), .S(n903) );
  CMPR32X2TF U1804 ( .A(b[6]), .B(b[7]), .C(n872), .CO(n871), .S(n904) );
  CMPR32X2TF U1805 ( .A(b[5]), .B(b[6]), .C(n873), .CO(n872), .S(n905) );
  CMPR32X2TF U1806 ( .A(b[4]), .B(b[5]), .C(n874), .CO(n873), .S(n906) );
  CMPR32X2TF U1807 ( .A(b[3]), .B(b[4]), .C(n875), .CO(n874), .S(n907) );
  CMPR32X2TF U1808 ( .A(b[2]), .B(b[3]), .C(n876), .CO(n875), .S(n908) );
  CMPR32X2TF U1809 ( .A(b[1]), .B(b[2]), .C(n877), .CO(n876), .S(n909) );
  ADDHXLTF U1810 ( .A(b[1]), .B(b[0]), .CO(n877), .S(n910) );
  OA21XLTF U1813 ( .A0(n2006), .A1(n127), .B0(n1292), .Y(n2289) );
  AOI22X1TF U1814 ( .A0(n3), .A1(n130), .B0(n1), .B1(n133), .Y(n2290) );
  AOI22X1TF U1815 ( .A0(n15), .A1(n130), .B0(n13), .B1(n133), .Y(n2291) );
  AOI22X1TF U1816 ( .A0(n27), .A1(n130), .B0(n25), .B1(n133), .Y(n2292) );
  AOI22X1TF U1817 ( .A0(n39), .A1(n130), .B0(n37), .B1(n133), .Y(n2293) );
  AOI22X1TF U1818 ( .A0(n51), .A1(n131), .B0(n49), .B1(n134), .Y(n2294) );
  AOI22X1TF U1819 ( .A0(n63), .A1(n131), .B0(n61), .B1(n134), .Y(n2295) );
  AOI22X1TF U1820 ( .A0(n75), .A1(n131), .B0(n73), .B1(n134), .Y(n2296) );
  AOI22X1TF U1821 ( .A0(n87), .A1(n132), .B0(n85), .B1(n134), .Y(n2297) );
  AOI22X1TF U1822 ( .A0(n99), .A1(n132), .B0(n97), .B1(n135), .Y(n2298) );
  AOI22X1TF U1823 ( .A0(n111), .A1(n132), .B0(n109), .B1(n135), .Y(n2299) );
  AOI22X1TF U1824 ( .A0(n123), .A1(n132), .B0(n121), .B1(n135), .Y(n2300) );
  NAND2X1TF U1825 ( .A(n1), .B(n130), .Y(n2301) );
  NAND2X1TF U1826 ( .A(n13), .B(n130), .Y(n2302) );
  NAND2X1TF U1827 ( .A(n25), .B(n130), .Y(n2303) );
  NAND2X1TF U1828 ( .A(n37), .B(n130), .Y(n2304) );
  NAND2X1TF U1829 ( .A(n49), .B(n131), .Y(n2305) );
  NAND2X1TF U1830 ( .A(n61), .B(n131), .Y(n2306) );
  NAND2X1TF U1831 ( .A(n73), .B(n131), .Y(n2307) );
  NAND2X1TF U1832 ( .A(n85), .B(n131), .Y(n2308) );
  NAND2X1TF U1833 ( .A(n97), .B(n132), .Y(n2309) );
  NAND2X1TF U1834 ( .A(n109), .B(n132), .Y(n2310) );
  NAND2X1TF U1835 ( .A(n121), .B(n132), .Y(n2311) );
  CLKBUFX2TF U1836 ( .A(n2147), .Y(n14) );
  CLKBUFX2TF U1837 ( .A(n2146), .Y(n26) );
  CLKBUFX2TF U1838 ( .A(n2145), .Y(n38) );
  CLKBUFX2TF U1839 ( .A(n2144), .Y(n50) );
  CLKBUFX2TF U1840 ( .A(n2143), .Y(n62) );
  CLKBUFX2TF U1841 ( .A(n2142), .Y(n74) );
  CLKBUFX2TF U1842 ( .A(n2141), .Y(n86) );
  CLKBUFX2TF U1843 ( .A(n2139), .Y(n110) );
  CLKBUFX2TF U1844 ( .A(n2140), .Y(n98) );
  CLKBUFX2TF U1845 ( .A(n2148), .Y(n2) );
  CLKBUFX2TF U1846 ( .A(n2146), .Y(n25) );
  CLKBUFX2TF U1847 ( .A(n2147), .Y(n13) );
  CLKBUFX2TF U1848 ( .A(n2144), .Y(n49) );
  CLKBUFX2TF U1849 ( .A(n2145), .Y(n37) );
  CLKBUFX2TF U1850 ( .A(n2142), .Y(n73) );
  CLKBUFX2TF U1851 ( .A(n2143), .Y(n61) );
  CLKBUFX2TF U1852 ( .A(n2140), .Y(n97) );
  CLKBUFX2TF U1853 ( .A(n2141), .Y(n85) );
  CLKBUFX2TF U1854 ( .A(n2139), .Y(n109) );
  CLKBUFX2TF U1855 ( .A(n2148), .Y(n1) );
  CLKBUFX2TF U1856 ( .A(n2124), .Y(n33) );
  CLKBUFX2TF U1857 ( .A(n2122), .Y(n57) );
  CLKBUFX2TF U1858 ( .A(n2125), .Y(n21) );
  CLKBUFX2TF U1859 ( .A(n2123), .Y(n45) );
  CLKBUFX2TF U1860 ( .A(n2121), .Y(n69) );
  CLKBUFX2TF U1861 ( .A(n2117), .Y(n117) );
  CLKBUFX2TF U1862 ( .A(n2118), .Y(n105) );
  CLKBUFX2TF U1863 ( .A(n2120), .Y(n81) );
  CLKBUFX2TF U1864 ( .A(n2119), .Y(n93) );
  CLKBUFX2TF U1865 ( .A(n2117), .Y(n118) );
  CLKBUFX2TF U1866 ( .A(n2125), .Y(n22) );
  CLKBUFX2TF U1867 ( .A(n2124), .Y(n34) );
  CLKBUFX2TF U1868 ( .A(n2123), .Y(n46) );
  CLKBUFX2TF U1869 ( .A(n2122), .Y(n58) );
  CLKBUFX2TF U1870 ( .A(n2121), .Y(n70) );
  CLKBUFX2TF U1871 ( .A(n2120), .Y(n82) );
  CLKBUFX2TF U1872 ( .A(n2119), .Y(n94) );
  CLKBUFX2TF U1873 ( .A(n2118), .Y(n106) );
  CLKBUFX2TF U1874 ( .A(n2126), .Y(n9) );
  CLKBUFX2TF U1875 ( .A(n2126), .Y(n10) );
  CLKBUFX2TF U1876 ( .A(n2136), .Y(n16) );
  CLKBUFX2TF U1877 ( .A(n2135), .Y(n28) );
  CLKBUFX2TF U1878 ( .A(n2134), .Y(n40) );
  CLKBUFX2TF U1879 ( .A(n2133), .Y(n52) );
  CLKBUFX2TF U1880 ( .A(n2132), .Y(n64) );
  CLKBUFX2TF U1881 ( .A(n2131), .Y(n76) );
  CLKBUFX2TF U1882 ( .A(n2130), .Y(n88) );
  CLKBUFX2TF U1883 ( .A(n2128), .Y(n112) );
  CLKBUFX2TF U1884 ( .A(n2129), .Y(n100) );
  CLKBUFX2TF U1885 ( .A(n2127), .Y(n124) );
  CLKBUFX2TF U1886 ( .A(n2137), .Y(n4) );
  CLKBUFX2TF U1887 ( .A(n2135), .Y(n27) );
  CLKBUFX2TF U1888 ( .A(n2136), .Y(n15) );
  CLKBUFX2TF U1889 ( .A(n2133), .Y(n51) );
  CLKBUFX2TF U1890 ( .A(n2134), .Y(n39) );
  CLKBUFX2TF U1891 ( .A(n2131), .Y(n75) );
  CLKBUFX2TF U1892 ( .A(n2132), .Y(n63) );
  CLKBUFX2TF U1893 ( .A(n2129), .Y(n99) );
  CLKBUFX2TF U1894 ( .A(n2130), .Y(n87) );
  CLKBUFX2TF U1895 ( .A(n2128), .Y(n111) );
  CLKBUFX2TF U1896 ( .A(n2127), .Y(n123) );
  CLKBUFX2TF U1897 ( .A(n2137), .Y(n3) );
  CLKBUFX2TF U1898 ( .A(n2124), .Y(n32) );
  CLKBUFX2TF U1899 ( .A(n2122), .Y(n56) );
  CLKBUFX2TF U1900 ( .A(n2125), .Y(n20) );
  CLKBUFX2TF U1901 ( .A(n2120), .Y(n80) );
  CLKBUFX2TF U1902 ( .A(n2123), .Y(n44) );
  CLKBUFX2TF U1903 ( .A(n2118), .Y(n104) );
  CLKBUFX2TF U1904 ( .A(n2121), .Y(n68) );
  CLKBUFX2TF U1905 ( .A(n2117), .Y(n116) );
  CLKBUFX2TF U1906 ( .A(n2119), .Y(n92) );
  CLKBUFX2TF U1907 ( .A(n2126), .Y(n8) );
  CLKBUFX2TF U1908 ( .A(n2113), .Y(n36) );
  CLKBUFX2TF U1909 ( .A(n2112), .Y(n48) );
  CLKBUFX2TF U1910 ( .A(n2111), .Y(n60) );
  CLKBUFX2TF U1911 ( .A(n2110), .Y(n72) );
  CLKBUFX2TF U1912 ( .A(n2109), .Y(n84) );
  CLKBUFX2TF U1913 ( .A(n2108), .Y(n96) );
  CLKBUFX2TF U1914 ( .A(n2106), .Y(n120) );
  CLKBUFX2TF U1915 ( .A(n2107), .Y(n108) );
  CLKBUFX2TF U1916 ( .A(n2114), .Y(n24) );
  CLKBUFX2TF U1917 ( .A(n2115), .Y(n12) );
  CLKBUFX2TF U1918 ( .A(n2113), .Y(n35) );
  CLKBUFX2TF U1919 ( .A(n2114), .Y(n23) );
  CLKBUFX2TF U1920 ( .A(n2111), .Y(n59) );
  CLKBUFX2TF U1921 ( .A(n2112), .Y(n47) );
  CLKBUFX2TF U1922 ( .A(n2109), .Y(n83) );
  CLKBUFX2TF U1923 ( .A(n2110), .Y(n71) );
  CLKBUFX2TF U1924 ( .A(n2107), .Y(n107) );
  CLKBUFX2TF U1925 ( .A(n2108), .Y(n95) );
  CLKBUFX2TF U1926 ( .A(n2106), .Y(n119) );
  CLKBUFX2TF U1927 ( .A(n2115), .Y(n11) );
  INVX2TF U1928 ( .A(n879), .Y(n2007) );
  INVX2TF U1929 ( .A(n910), .Y(n2038) );
  INVX2TF U1930 ( .A(n878), .Y(n2006) );
  INVX2TF U1931 ( .A(n909), .Y(n2037) );
  INVX2TF U1932 ( .A(n908), .Y(n2036) );
  INVX2TF U1933 ( .A(n907), .Y(n2035) );
  INVX2TF U1934 ( .A(n906), .Y(n2034) );
  INVX2TF U1935 ( .A(n905), .Y(n2033) );
  INVX2TF U1936 ( .A(n903), .Y(n2031) );
  INVX2TF U1937 ( .A(n904), .Y(n2032) );
  INVX2TF U1938 ( .A(n898), .Y(n2026) );
  INVX2TF U1939 ( .A(n897), .Y(n2025) );
  INVX2TF U1940 ( .A(n902), .Y(n2030) );
  INVX2TF U1941 ( .A(n901), .Y(n2029) );
  INVX2TF U1942 ( .A(n900), .Y(n2028) );
  INVX2TF U1943 ( .A(n899), .Y(n2027) );
  INVX2TF U1944 ( .A(n892), .Y(n2020) );
  INVX2TF U1945 ( .A(n891), .Y(n2019) );
  INVX2TF U1946 ( .A(n895), .Y(n2023) );
  INVX2TF U1947 ( .A(n894), .Y(n2022) );
  INVX2TF U1948 ( .A(n896), .Y(n2024) );
  INVX2TF U1949 ( .A(n893), .Y(n2021) );
  INVX2TF U1950 ( .A(n888), .Y(n2016) );
  INVX2TF U1951 ( .A(n890), .Y(n2018) );
  INVX2TF U1952 ( .A(n889), .Y(n2017) );
  INVX2TF U1953 ( .A(n887), .Y(n2015) );
  INVX2TF U1954 ( .A(n886), .Y(n2014) );
  INVX2TF U1955 ( .A(n880), .Y(n2008) );
  INVX2TF U1956 ( .A(n885), .Y(n2013) );
  INVX2TF U1957 ( .A(n884), .Y(n2012) );
  INVX2TF U1958 ( .A(n883), .Y(n2011) );
  INVX2TF U1959 ( .A(n882), .Y(n2010) );
  INVX2TF U1960 ( .A(n881), .Y(n2009) );
  CLKBUFX2TF U1961 ( .A(n2138), .Y(n122) );
  CLKBUFX2TF U1962 ( .A(n2138), .Y(n121) );
  CLKBUFX2TF U1963 ( .A(n2116), .Y(n126) );
  CLKBUFX2TF U1964 ( .A(n2116), .Y(n127) );
  CLKBUFX2TF U1965 ( .A(n2116), .Y(n125) );
  CLKBUFX2TF U1966 ( .A(n2158), .Y(n7) );
  CLKBUFX2TF U1967 ( .A(n2105), .Y(n129) );
  CLKBUFX2TF U1968 ( .A(n2105), .Y(n128) );
  CLKBUFX2TF U1969 ( .A(n2158), .Y(n5) );
  CLKBUFX2TF U1970 ( .A(n2158), .Y(n6) );
  CLKBUFX2TF U1971 ( .A(n2157), .Y(n19) );
  CLKBUFX2TF U1972 ( .A(n2156), .Y(n31) );
  CLKBUFX2TF U1973 ( .A(n2155), .Y(n43) );
  CLKBUFX2TF U1974 ( .A(n2154), .Y(n55) );
  CLKBUFX2TF U1975 ( .A(n2153), .Y(n67) );
  CLKBUFX2TF U1976 ( .A(n2152), .Y(n79) );
  CLKBUFX2TF U1977 ( .A(n2151), .Y(n91) );
  CLKBUFX2TF U1978 ( .A(n2150), .Y(n103) );
  CLKBUFX2TF U1979 ( .A(n2149), .Y(n115) );
  CLKBUFX2TF U1980 ( .A(n2157), .Y(n17) );
  CLKBUFX2TF U1981 ( .A(n2155), .Y(n41) );
  CLKBUFX2TF U1982 ( .A(n2153), .Y(n65) );
  CLKBUFX2TF U1983 ( .A(n2157), .Y(n18) );
  CLKBUFX2TF U1984 ( .A(n2156), .Y(n29) );
  CLKBUFX2TF U1985 ( .A(n2151), .Y(n89) );
  CLKBUFX2TF U1986 ( .A(n2155), .Y(n42) );
  CLKBUFX2TF U1987 ( .A(n2154), .Y(n53) );
  CLKBUFX2TF U1988 ( .A(n2152), .Y(n77) );
  CLKBUFX2TF U1989 ( .A(n2150), .Y(n101) );
  CLKBUFX2TF U1990 ( .A(n2156), .Y(n30) );
  CLKBUFX2TF U1991 ( .A(n2149), .Y(n113) );
  CLKBUFX2TF U1992 ( .A(n2154), .Y(n54) );
  CLKBUFX2TF U1993 ( .A(n2153), .Y(n66) );
  CLKBUFX2TF U1994 ( .A(n2152), .Y(n78) );
  CLKBUFX2TF U1995 ( .A(n2151), .Y(n90) );
  CLKBUFX2TF U1996 ( .A(n2150), .Y(n102) );
  CLKBUFX2TF U1997 ( .A(n2149), .Y(n114) );
  CLKBUFX2TF U1998 ( .A(n2040), .Y(n225) );
  CLKBUFX2TF U1999 ( .A(n2040), .Y(n224) );
  CLKBUFX2TF U2000 ( .A(n2041), .Y(n221) );
  CLKBUFX2TF U2001 ( .A(n2041), .Y(n222) );
  CLKBUFX2TF U2002 ( .A(n2040), .Y(n223) );
  CLKBUFX2TF U2003 ( .A(n2041), .Y(n220) );
  CLKBUFX2TF U2004 ( .A(n2069), .Y(n136) );
  CLKBUFX2TF U2005 ( .A(n2068), .Y(n139) );
  CLKBUFX2TF U2006 ( .A(n2067), .Y(n142) );
  CLKBUFX2TF U2007 ( .A(n2066), .Y(n145) );
  CLKBUFX2TF U2008 ( .A(n2065), .Y(n148) );
  CLKBUFX2TF U2009 ( .A(n2064), .Y(n151) );
  CLKBUFX2TF U2010 ( .A(n2063), .Y(n154) );
  CLKBUFX2TF U2011 ( .A(n2062), .Y(n157) );
  CLKBUFX2TF U2012 ( .A(n2061), .Y(n160) );
  CLKBUFX2TF U2013 ( .A(n2060), .Y(n163) );
  CLKBUFX2TF U2014 ( .A(n2059), .Y(n166) );
  CLKBUFX2TF U2015 ( .A(n2058), .Y(n169) );
  CLKBUFX2TF U2016 ( .A(n2057), .Y(n172) );
  CLKBUFX2TF U2017 ( .A(n2056), .Y(n175) );
  CLKBUFX2TF U2018 ( .A(n2055), .Y(n178) );
  CLKBUFX2TF U2019 ( .A(n2054), .Y(n181) );
  CLKBUFX2TF U2020 ( .A(n2053), .Y(n184) );
  CLKBUFX2TF U2021 ( .A(n2052), .Y(n187) );
  CLKBUFX2TF U2022 ( .A(n2051), .Y(n190) );
  CLKBUFX2TF U2023 ( .A(n2050), .Y(n193) );
  CLKBUFX2TF U2024 ( .A(n2049), .Y(n196) );
  CLKBUFX2TF U2025 ( .A(n2048), .Y(n199) );
  CLKBUFX2TF U2026 ( .A(n2047), .Y(n202) );
  CLKBUFX2TF U2027 ( .A(n2046), .Y(n205) );
  CLKBUFX2TF U2028 ( .A(n2045), .Y(n208) );
  CLKBUFX2TF U2029 ( .A(n2044), .Y(n211) );
  CLKBUFX2TF U2030 ( .A(n2043), .Y(n214) );
  CLKBUFX2TF U2031 ( .A(n2042), .Y(n217) );
  CLKBUFX2TF U2032 ( .A(n2065), .Y(n149) );
  CLKBUFX2TF U2033 ( .A(n2064), .Y(n152) );
  CLKBUFX2TF U2034 ( .A(n2063), .Y(n155) );
  CLKBUFX2TF U2035 ( .A(n2062), .Y(n158) );
  CLKBUFX2TF U2036 ( .A(n2069), .Y(n137) );
  CLKBUFX2TF U2037 ( .A(n2061), .Y(n161) );
  CLKBUFX2TF U2038 ( .A(n2068), .Y(n140) );
  CLKBUFX2TF U2039 ( .A(n2060), .Y(n164) );
  CLKBUFX2TF U2040 ( .A(n2067), .Y(n143) );
  CLKBUFX2TF U2041 ( .A(n2059), .Y(n167) );
  CLKBUFX2TF U2042 ( .A(n2066), .Y(n146) );
  CLKBUFX2TF U2043 ( .A(n2058), .Y(n170) );
  CLKBUFX2TF U2044 ( .A(n2057), .Y(n173) );
  CLKBUFX2TF U2045 ( .A(n2056), .Y(n176) );
  CLKBUFX2TF U2046 ( .A(n2055), .Y(n179) );
  CLKBUFX2TF U2047 ( .A(n2054), .Y(n182) );
  CLKBUFX2TF U2048 ( .A(n2053), .Y(n185) );
  CLKBUFX2TF U2049 ( .A(n2052), .Y(n188) );
  CLKBUFX2TF U2050 ( .A(n2051), .Y(n191) );
  CLKBUFX2TF U2051 ( .A(n2050), .Y(n194) );
  CLKBUFX2TF U2052 ( .A(n2048), .Y(n200) );
  CLKBUFX2TF U2053 ( .A(n2049), .Y(n197) );
  CLKBUFX2TF U2054 ( .A(n2047), .Y(n203) );
  CLKBUFX2TF U2055 ( .A(n2046), .Y(n206) );
  CLKBUFX2TF U2056 ( .A(n2045), .Y(n209) );
  CLKBUFX2TF U2057 ( .A(n2044), .Y(n212) );
  CLKBUFX2TF U2058 ( .A(n2043), .Y(n215) );
  CLKBUFX2TF U2059 ( .A(n2042), .Y(n218) );
  CLKBUFX2TF U2060 ( .A(n2066), .Y(n147) );
  CLKBUFX2TF U2061 ( .A(n2065), .Y(n150) );
  CLKBUFX2TF U2062 ( .A(n2064), .Y(n153) );
  CLKBUFX2TF U2063 ( .A(n2063), .Y(n156) );
  CLKBUFX2TF U2064 ( .A(n2062), .Y(n159) );
  CLKBUFX2TF U2065 ( .A(n2061), .Y(n162) );
  CLKBUFX2TF U2066 ( .A(n2069), .Y(n138) );
  CLKBUFX2TF U2067 ( .A(n2068), .Y(n141) );
  CLKBUFX2TF U2068 ( .A(n2067), .Y(n144) );
  CLKBUFX2TF U2069 ( .A(n2056), .Y(n177) );
  CLKBUFX2TF U2070 ( .A(n2060), .Y(n165) );
  CLKBUFX2TF U2071 ( .A(n2059), .Y(n168) );
  CLKBUFX2TF U2072 ( .A(n2058), .Y(n171) );
  CLKBUFX2TF U2073 ( .A(n2055), .Y(n180) );
  CLKBUFX2TF U2074 ( .A(n2057), .Y(n174) );
  CLKBUFX2TF U2075 ( .A(n2054), .Y(n183) );
  CLKBUFX2TF U2076 ( .A(n2053), .Y(n186) );
  CLKBUFX2TF U2077 ( .A(n2052), .Y(n189) );
  CLKBUFX2TF U2078 ( .A(n2051), .Y(n192) );
  CLKBUFX2TF U2079 ( .A(n2050), .Y(n195) );
  CLKBUFX2TF U2080 ( .A(n2045), .Y(n210) );
  CLKBUFX2TF U2081 ( .A(n2046), .Y(n207) );
  CLKBUFX2TF U2082 ( .A(n2049), .Y(n198) );
  CLKBUFX2TF U2083 ( .A(n2048), .Y(n201) );
  CLKBUFX2TF U2084 ( .A(n2047), .Y(n204) );
  CLKBUFX2TF U2085 ( .A(n2044), .Y(n213) );
  CLKBUFX2TF U2086 ( .A(n2043), .Y(n216) );
  CLKBUFX2TF U2087 ( .A(n2042), .Y(n219) );
  CLKBUFX2TF U2088 ( .A(n2071), .Y(n131) );
  CLKBUFX2TF U2089 ( .A(n2071), .Y(n130) );
  CLKBUFX2TF U2090 ( .A(n2071), .Y(n132) );
  CLKBUFX2TF U2091 ( .A(n2070), .Y(n135) );
  CLKBUFX2TF U2092 ( .A(n2070), .Y(n133) );
  CLKBUFX2TF U2093 ( .A(n2070), .Y(n134) );
  CLKBUFX2TF U2094 ( .A(a[5]), .Y(n2157) );
  CLKBUFX2TF U2095 ( .A(a[11]), .Y(n2155) );
  CLKBUFX2TF U2096 ( .A(a[17]), .Y(n2153) );
  CLKBUFX2TF U2097 ( .A(a[8]), .Y(n2156) );
  CLKBUFX2TF U2098 ( .A(a[23]), .Y(n2151) );
  CLKBUFX2TF U2099 ( .A(b[5]), .Y(n2066) );
  CLKBUFX2TF U2100 ( .A(a[14]), .Y(n2154) );
  CLKBUFX2TF U2101 ( .A(b[6]), .Y(n2065) );
  CLKBUFX2TF U2102 ( .A(b[7]), .Y(n2064) );
  CLKBUFX2TF U2103 ( .A(b[8]), .Y(n2063) );
  CLKBUFX2TF U2104 ( .A(b[9]), .Y(n2062) );
  CLKBUFX2TF U2105 ( .A(b[0]), .Y(n2071) );
  CLKBUFX2TF U2106 ( .A(a[20]), .Y(n2152) );
  CLKBUFX2TF U2107 ( .A(b[10]), .Y(n2061) );
  CLKBUFX2TF U2108 ( .A(b[1]), .Y(n2070) );
  CLKBUFX2TF U2109 ( .A(b[2]), .Y(n2069) );
  CLKBUFX2TF U2110 ( .A(b[3]), .Y(n2068) );
  CLKBUFX2TF U2111 ( .A(b[4]), .Y(n2067) );
  CLKBUFX2TF U2112 ( .A(a[26]), .Y(n2150) );
  CLKBUFX2TF U2113 ( .A(b[15]), .Y(n2056) );
  CLKBUFX2TF U2114 ( .A(b[11]), .Y(n2060) );
  CLKBUFX2TF U2115 ( .A(b[12]), .Y(n2059) );
  CLKBUFX2TF U2116 ( .A(b[13]), .Y(n2058) );
  CLKBUFX2TF U2117 ( .A(a[29]), .Y(n2149) );
  CLKBUFX2TF U2118 ( .A(b[16]), .Y(n2055) );
  CLKBUFX2TF U2119 ( .A(b[14]), .Y(n2057) );
  CLKBUFX2TF U2120 ( .A(b[17]), .Y(n2054) );
  CLKBUFX2TF U2121 ( .A(b[18]), .Y(n2053) );
  CLKBUFX2TF U2122 ( .A(b[19]), .Y(n2052) );
  CLKBUFX2TF U2123 ( .A(b[20]), .Y(n2051) );
  CLKBUFX2TF U2124 ( .A(b[21]), .Y(n2050) );
  CLKBUFX2TF U2125 ( .A(b[26]), .Y(n2045) );
  CLKBUFX2TF U2126 ( .A(b[25]), .Y(n2046) );
  CLKBUFX2TF U2127 ( .A(b[22]), .Y(n2049) );
  CLKBUFX2TF U2128 ( .A(b[23]), .Y(n2048) );
  CLKBUFX2TF U2129 ( .A(b[24]), .Y(n2047) );
  CLKBUFX2TF U2130 ( .A(b[27]), .Y(n2044) );
  CLKBUFX2TF U2131 ( .A(b[28]), .Y(n2043) );
  CLKBUFX2TF U2132 ( .A(b[31]), .Y(n2040) );
  CLKBUFX2TF U2133 ( .A(b[30]), .Y(n2041) );
  CLKBUFX2TF U2134 ( .A(b[29]), .Y(n2042) );
  CLKBUFX2TF U2135 ( .A(a[2]), .Y(n2158) );
  INVX2TF U2136 ( .A(b[0]), .Y(n2039) );
endmodule


module mul ( A, B, X );
  input [31:0] A;
  input [31:0] B;
  output [63:0] X;


  mul_DW_mult_uns_1 mult_3 ( .a(A), .b(B), .product(X) );
endmodule

