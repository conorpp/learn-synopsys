module mul(input[31:0] A,input[31:0] B, output[63:0] X);

assign X = A * B;

endmodule
